module rom(
    input i_clk_a,
    input[14:0] i_addr_a,
    output reg[15:0] o_data_a
);

   always @* begin
       case (i_addr_a)
            14'h0000: o_data_a = 16'b0000000100000000;
            14'h0001: o_data_a = 16'b1110110000010000;
            14'h0002: o_data_a = 16'b0000000000000000;
            14'h0003: o_data_a = 16'b1110001100001000;
            14'h0004: o_data_a = 16'b0000000010000101;
            14'h0005: o_data_a = 16'b1110101010000111;
            14'h0006: o_data_a = 16'b0000000000001111;
            14'h0007: o_data_a = 16'b1110001100001000;
            14'h0008: o_data_a = 16'b0000000000000000;
            14'h0009: o_data_a = 16'b1111110010101000;
            14'h000a: o_data_a = 16'b1111110000010000;
            14'h000b: o_data_a = 16'b1110110010100000;
            14'h000c: o_data_a = 16'b1111000111010000;
            14'h000d: o_data_a = 16'b1110101010001000;
            14'h000e: o_data_a = 16'b0000000000010011;
            14'h000f: o_data_a = 16'b1110001100000101;
            14'h0010: o_data_a = 16'b0000000000000000;
            14'h0011: o_data_a = 16'b1111110010100000;
            14'h0012: o_data_a = 16'b1110111010001000;
            14'h0013: o_data_a = 16'b0000000000001111;
            14'h0014: o_data_a = 16'b1111110000100000;
            14'h0015: o_data_a = 16'b1110101010000111;
            14'h0016: o_data_a = 16'b0000000000001111;
            14'h0017: o_data_a = 16'b1110001100001000;
            14'h0018: o_data_a = 16'b0000000000000000;
            14'h0019: o_data_a = 16'b1111110010101000;
            14'h001a: o_data_a = 16'b1111110000010000;
            14'h001b: o_data_a = 16'b1110110010100000;
            14'h001c: o_data_a = 16'b1111000111010000;
            14'h001d: o_data_a = 16'b1110101010001000;
            14'h001e: o_data_a = 16'b0000000000100011;
            14'h001f: o_data_a = 16'b1110001100000110;
            14'h0020: o_data_a = 16'b0000000000000000;
            14'h0021: o_data_a = 16'b1111110010100000;
            14'h0022: o_data_a = 16'b1110111010001000;
            14'h0023: o_data_a = 16'b0000000000001111;
            14'h0024: o_data_a = 16'b1111110000100000;
            14'h0025: o_data_a = 16'b1110101010000111;
            14'h0026: o_data_a = 16'b0000000000001111;
            14'h0027: o_data_a = 16'b1110001100001000;
            14'h0028: o_data_a = 16'b0000000000000000;
            14'h0029: o_data_a = 16'b1111110010101000;
            14'h002a: o_data_a = 16'b1111110000010000;
            14'h002b: o_data_a = 16'b1110110010100000;
            14'h002c: o_data_a = 16'b1111000111010000;
            14'h002d: o_data_a = 16'b1110101010001000;
            14'h002e: o_data_a = 16'b0000000000110011;
            14'h002f: o_data_a = 16'b1110001100000011;
            14'h0030: o_data_a = 16'b0000000000000000;
            14'h0031: o_data_a = 16'b1111110010100000;
            14'h0032: o_data_a = 16'b1110111010001000;
            14'h0033: o_data_a = 16'b0000000000001111;
            14'h0034: o_data_a = 16'b1111110000100000;
            14'h0035: o_data_a = 16'b1110101010000111;
            14'h0036: o_data_a = 16'b0000000000000101;
            14'h0037: o_data_a = 16'b1110110000010000;
            14'h0038: o_data_a = 16'b0000000000000001;
            14'h0039: o_data_a = 16'b1111000111100000;
            14'h003a: o_data_a = 16'b1111110000010000;
            14'h003b: o_data_a = 16'b0000000000001101;
            14'h003c: o_data_a = 16'b1110001100001000;
            14'h003d: o_data_a = 16'b0000000000000000;
            14'h003e: o_data_a = 16'b1111110010101000;
            14'h003f: o_data_a = 16'b1111110000010000;
            14'h0040: o_data_a = 16'b0000000000000010;
            14'h0041: o_data_a = 16'b1111110000100000;
            14'h0042: o_data_a = 16'b1110001100001000;
            14'h0043: o_data_a = 16'b1110110000010000;
            14'h0044: o_data_a = 16'b0000000000000000;
            14'h0045: o_data_a = 16'b1110011111001000;
            14'h0046: o_data_a = 16'b0000000000000001;
            14'h0047: o_data_a = 16'b1111110000010000;
            14'h0048: o_data_a = 16'b0000000000001110;
            14'h0049: o_data_a = 16'b1110001110101000;
            14'h004a: o_data_a = 16'b1111110000010000;
            14'h004b: o_data_a = 16'b0000000000000100;
            14'h004c: o_data_a = 16'b1110001100001000;
            14'h004d: o_data_a = 16'b0000000000001110;
            14'h004e: o_data_a = 16'b1111110010101000;
            14'h004f: o_data_a = 16'b1111110000010000;
            14'h0050: o_data_a = 16'b0000000000000011;
            14'h0051: o_data_a = 16'b1110001100001000;
            14'h0052: o_data_a = 16'b0000000000001110;
            14'h0053: o_data_a = 16'b1111110010101000;
            14'h0054: o_data_a = 16'b1111110000010000;
            14'h0055: o_data_a = 16'b0000000000000010;
            14'h0056: o_data_a = 16'b1110001100001000;
            14'h0057: o_data_a = 16'b0000000000001110;
            14'h0058: o_data_a = 16'b1111110010101000;
            14'h0059: o_data_a = 16'b1111110000010000;
            14'h005a: o_data_a = 16'b0000000000000001;
            14'h005b: o_data_a = 16'b1110001100001000;
            14'h005c: o_data_a = 16'b0000000000001101;
            14'h005d: o_data_a = 16'b1111110000100000;
            14'h005e: o_data_a = 16'b1110101010000111;
            14'h005f: o_data_a = 16'b0000000000000000;
            14'h0060: o_data_a = 16'b1111110000100000;
            14'h0061: o_data_a = 16'b1110001100001000;
            14'h0062: o_data_a = 16'b0000000000000001;
            14'h0063: o_data_a = 16'b1111110000010000;
            14'h0064: o_data_a = 16'b0000000000000000;
            14'h0065: o_data_a = 16'b1111110111101000;
            14'h0066: o_data_a = 16'b1110001100001000;
            14'h0067: o_data_a = 16'b0000000000000010;
            14'h0068: o_data_a = 16'b1111110000010000;
            14'h0069: o_data_a = 16'b0000000000000000;
            14'h006a: o_data_a = 16'b1111110111101000;
            14'h006b: o_data_a = 16'b1110001100001000;
            14'h006c: o_data_a = 16'b0000000000000011;
            14'h006d: o_data_a = 16'b1111110000010000;
            14'h006e: o_data_a = 16'b0000000000000000;
            14'h006f: o_data_a = 16'b1111110111101000;
            14'h0070: o_data_a = 16'b1110001100001000;
            14'h0071: o_data_a = 16'b0000000000000100;
            14'h0072: o_data_a = 16'b1111110000010000;
            14'h0073: o_data_a = 16'b0000000000000000;
            14'h0074: o_data_a = 16'b1111110111101000;
            14'h0075: o_data_a = 16'b1110001100001000;
            14'h0076: o_data_a = 16'b0000000000000100;
            14'h0077: o_data_a = 16'b1110110000010000;
            14'h0078: o_data_a = 16'b0000000000001101;
            14'h0079: o_data_a = 16'b1111000010010000;
            14'h007a: o_data_a = 16'b0000000000000000;
            14'h007b: o_data_a = 16'b1111000111010000;
            14'h007c: o_data_a = 16'b0000000000000010;
            14'h007d: o_data_a = 16'b1110001100001000;
            14'h007e: o_data_a = 16'b0000000000000000;
            14'h007f: o_data_a = 16'b1111110111011000;
            14'h0080: o_data_a = 16'b0000000000000001;
            14'h0081: o_data_a = 16'b1110001100001000;
            14'h0082: o_data_a = 16'b0000000000001110;
            14'h0083: o_data_a = 16'b1111110000100000;
            14'h0084: o_data_a = 16'b1110101010000111;
            14'h0085: o_data_a = 16'b0000000000000000;
            14'h0086: o_data_a = 16'b1110110000010000;
            14'h0087: o_data_a = 16'b0000000000001101;
            14'h0088: o_data_a = 16'b1110001100001000;
            14'h0089: o_data_a = 16'b0110100110110010;
            14'h008a: o_data_a = 16'b1110110000010000;
            14'h008b: o_data_a = 16'b0000000000001110;
            14'h008c: o_data_a = 16'b1110001100001000;
            14'h008d: o_data_a = 16'b0000000010010001;
            14'h008e: o_data_a = 16'b1110110000010000;
            14'h008f: o_data_a = 16'b0000000001011111;
            14'h0090: o_data_a = 16'b1110101010000111;
            14'h0091: o_data_a = 16'b0000000000001111;
            14'h0092: o_data_a = 16'b1110110000010000;
            14'h0093: o_data_a = 16'b0000000000000000;
            14'h0094: o_data_a = 16'b1111110111101000;
            14'h0095: o_data_a = 16'b1110110010100000;
            14'h0096: o_data_a = 16'b1110001100001000;
            14'h0097: o_data_a = 16'b0000000000000001;
            14'h0098: o_data_a = 16'b1110110000010000;
            14'h0099: o_data_a = 16'b0000000000001101;
            14'h009a: o_data_a = 16'b1110001100001000;
            14'h009b: o_data_a = 16'b0010000111000011;
            14'h009c: o_data_a = 16'b1110110000010000;
            14'h009d: o_data_a = 16'b0000000000001110;
            14'h009e: o_data_a = 16'b1110001100001000;
            14'h009f: o_data_a = 16'b0000000010100011;
            14'h00a0: o_data_a = 16'b1110110000010000;
            14'h00a1: o_data_a = 16'b0000000001011111;
            14'h00a2: o_data_a = 16'b1110101010000111;
            14'h00a3: o_data_a = 16'b0000000000000000;
            14'h00a4: o_data_a = 16'b1111110010101000;
            14'h00a5: o_data_a = 16'b1111110000010000;
            14'h00a6: o_data_a = 16'b0000000000000011;
            14'h00a7: o_data_a = 16'b1110001100001000;
            14'h00a8: o_data_a = 16'b0000000000000010;
            14'h00a9: o_data_a = 16'b1111110000100000;
            14'h00aa: o_data_a = 16'b1111110000010000;
            14'h00ab: o_data_a = 16'b0000000000000000;
            14'h00ac: o_data_a = 16'b1111110111101000;
            14'h00ad: o_data_a = 16'b1110110010100000;
            14'h00ae: o_data_a = 16'b1110001100001000;
            14'h00af: o_data_a = 16'b0000000000000000;
            14'h00b0: o_data_a = 16'b1111110010101000;
            14'h00b1: o_data_a = 16'b1111110000010000;
            14'h00b2: o_data_a = 16'b0000000000000011;
            14'h00b3: o_data_a = 16'b1111110000100000;
            14'h00b4: o_data_a = 16'b1110001100001000;
            14'h00b5: o_data_a = 16'b0000000000000010;
            14'h00b6: o_data_a = 16'b1111110111100000;
            14'h00b7: o_data_a = 16'b1111110000010000;
            14'h00b8: o_data_a = 16'b0000000000000000;
            14'h00b9: o_data_a = 16'b1111110111101000;
            14'h00ba: o_data_a = 16'b1110110010100000;
            14'h00bb: o_data_a = 16'b1110001100001000;
            14'h00bc: o_data_a = 16'b0000000000000000;
            14'h00bd: o_data_a = 16'b1111110010101000;
            14'h00be: o_data_a = 16'b1111110000010000;
            14'h00bf: o_data_a = 16'b0000000000000011;
            14'h00c0: o_data_a = 16'b1111110111100000;
            14'h00c1: o_data_a = 16'b1110001100001000;
            14'h00c2: o_data_a = 16'b0000000000000010;
            14'h00c3: o_data_a = 16'b1111110111100000;
            14'h00c4: o_data_a = 16'b1110110111100000;
            14'h00c5: o_data_a = 16'b1111110000010000;
            14'h00c6: o_data_a = 16'b0000000000000000;
            14'h00c7: o_data_a = 16'b1111110111101000;
            14'h00c8: o_data_a = 16'b1110110010100000;
            14'h00c9: o_data_a = 16'b1110001100001000;
            14'h00ca: o_data_a = 16'b0000000000000011;
            14'h00cb: o_data_a = 16'b1111110000010000;
            14'h00cc: o_data_a = 16'b0000000000001010;
            14'h00cd: o_data_a = 16'b1110000010010000;
            14'h00ce: o_data_a = 16'b0000000000001101;
            14'h00cf: o_data_a = 16'b1110001100001000;
            14'h00d0: o_data_a = 16'b0000000000000000;
            14'h00d1: o_data_a = 16'b1111110010101000;
            14'h00d2: o_data_a = 16'b1111110000010000;
            14'h00d3: o_data_a = 16'b0000000000001101;
            14'h00d4: o_data_a = 16'b1111110000100000;
            14'h00d5: o_data_a = 16'b1110001100001000;
            14'h00d6: o_data_a = 16'b0000000000000010;
            14'h00d7: o_data_a = 16'b1111110000010000;
            14'h00d8: o_data_a = 16'b0000000000000011;
            14'h00d9: o_data_a = 16'b1110000010100000;
            14'h00da: o_data_a = 16'b1111110000010000;
            14'h00db: o_data_a = 16'b0000000000000000;
            14'h00dc: o_data_a = 16'b1111110111101000;
            14'h00dd: o_data_a = 16'b1110110010100000;
            14'h00de: o_data_a = 16'b1110001100001000;
            14'h00df: o_data_a = 16'b0000000000000110;
            14'h00e0: o_data_a = 16'b1110110000010000;
            14'h00e1: o_data_a = 16'b0000000000000000;
            14'h00e2: o_data_a = 16'b1111110111101000;
            14'h00e3: o_data_a = 16'b1110110010100000;
            14'h00e4: o_data_a = 16'b1110001100001000;
            14'h00e5: o_data_a = 16'b0000000000000000;
            14'h00e6: o_data_a = 16'b1111110010101000;
            14'h00e7: o_data_a = 16'b1111110000010000;
            14'h00e8: o_data_a = 16'b1110110010100000;
            14'h00e9: o_data_a = 16'b1111000111001000;
            14'h00ea: o_data_a = 16'b0000000000000011;
            14'h00eb: o_data_a = 16'b1111110000010000;
            14'h00ec: o_data_a = 16'b0000000000001011;
            14'h00ed: o_data_a = 16'b1110000010010000;
            14'h00ee: o_data_a = 16'b0000000000001101;
            14'h00ef: o_data_a = 16'b1110001100001000;
            14'h00f0: o_data_a = 16'b0000000000000000;
            14'h00f1: o_data_a = 16'b1111110010101000;
            14'h00f2: o_data_a = 16'b1111110000010000;
            14'h00f3: o_data_a = 16'b0000000000001101;
            14'h00f4: o_data_a = 16'b1111110000100000;
            14'h00f5: o_data_a = 16'b1110001100001000;
            14'h00f6: o_data_a = 16'b0000000000000010;
            14'h00f7: o_data_a = 16'b1111110000010000;
            14'h00f8: o_data_a = 16'b0000000000000100;
            14'h00f9: o_data_a = 16'b1110000010100000;
            14'h00fa: o_data_a = 16'b1111110000010000;
            14'h00fb: o_data_a = 16'b0000000000000000;
            14'h00fc: o_data_a = 16'b1111110111101000;
            14'h00fd: o_data_a = 16'b1110110010100000;
            14'h00fe: o_data_a = 16'b1110001100001000;
            14'h00ff: o_data_a = 16'b0000000000000011;
            14'h0100: o_data_a = 16'b1111110000010000;
            14'h0101: o_data_a = 16'b0000000000001100;
            14'h0102: o_data_a = 16'b1110000010010000;
            14'h0103: o_data_a = 16'b0000000000001101;
            14'h0104: o_data_a = 16'b1110001100001000;
            14'h0105: o_data_a = 16'b0000000000000000;
            14'h0106: o_data_a = 16'b1111110010101000;
            14'h0107: o_data_a = 16'b1111110000010000;
            14'h0108: o_data_a = 16'b0000000000001101;
            14'h0109: o_data_a = 16'b1111110000100000;
            14'h010a: o_data_a = 16'b1110001100001000;
            14'h010b: o_data_a = 16'b0000000000000010;
            14'h010c: o_data_a = 16'b1111110000010000;
            14'h010d: o_data_a = 16'b0000000000000101;
            14'h010e: o_data_a = 16'b1110000010100000;
            14'h010f: o_data_a = 16'b1111110000010000;
            14'h0110: o_data_a = 16'b0000000000000000;
            14'h0111: o_data_a = 16'b1111110111101000;
            14'h0112: o_data_a = 16'b1110110010100000;
            14'h0113: o_data_a = 16'b1110001100001000;
            14'h0114: o_data_a = 16'b0000000000000110;
            14'h0115: o_data_a = 16'b1110110000010000;
            14'h0116: o_data_a = 16'b0000000000000000;
            14'h0117: o_data_a = 16'b1111110111101000;
            14'h0118: o_data_a = 16'b1110110010100000;
            14'h0119: o_data_a = 16'b1110001100001000;
            14'h011a: o_data_a = 16'b0000000000000000;
            14'h011b: o_data_a = 16'b1111110010101000;
            14'h011c: o_data_a = 16'b1111110000010000;
            14'h011d: o_data_a = 16'b1110110010100000;
            14'h011e: o_data_a = 16'b1111000111001000;
            14'h011f: o_data_a = 16'b0000000000000011;
            14'h0120: o_data_a = 16'b1111110000010000;
            14'h0121: o_data_a = 16'b0000000000001101;
            14'h0122: o_data_a = 16'b1110000010010000;
            14'h0123: o_data_a = 16'b0000000000001101;
            14'h0124: o_data_a = 16'b1110001100001000;
            14'h0125: o_data_a = 16'b0000000000000000;
            14'h0126: o_data_a = 16'b1111110010101000;
            14'h0127: o_data_a = 16'b1111110000010000;
            14'h0128: o_data_a = 16'b0000000000001101;
            14'h0129: o_data_a = 16'b1111110000100000;
            14'h012a: o_data_a = 16'b1110001100001000;
            14'h012b: o_data_a = 16'b0000000000000000;
            14'h012c: o_data_a = 16'b1111110111001000;
            14'h012d: o_data_a = 16'b1111110010100000;
            14'h012e: o_data_a = 16'b1110101010001000;
            14'h012f: o_data_a = 16'b0000000000000011;
            14'h0130: o_data_a = 16'b1111110000010000;
            14'h0131: o_data_a = 16'b0000000000001110;
            14'h0132: o_data_a = 16'b1110000010010000;
            14'h0133: o_data_a = 16'b0000000000001101;
            14'h0134: o_data_a = 16'b1110001100001000;
            14'h0135: o_data_a = 16'b0000000000000000;
            14'h0136: o_data_a = 16'b1111110010101000;
            14'h0137: o_data_a = 16'b1111110000010000;
            14'h0138: o_data_a = 16'b0000000000001101;
            14'h0139: o_data_a = 16'b1111110000100000;
            14'h013a: o_data_a = 16'b1110001100001000;
            14'h013b: o_data_a = 16'b0000000000000011;
            14'h013c: o_data_a = 16'b1111110000010000;
            14'h013d: o_data_a = 16'b0000000000000000;
            14'h013e: o_data_a = 16'b1111110111101000;
            14'h013f: o_data_a = 16'b1110110010100000;
            14'h0140: o_data_a = 16'b1110001100001000;
            14'h0141: o_data_a = 16'b0000000000000001;
            14'h0142: o_data_a = 16'b1110110000010000;
            14'h0143: o_data_a = 16'b0000000000001101;
            14'h0144: o_data_a = 16'b1110001100001000;
            14'h0145: o_data_a = 16'b0000000110000011;
            14'h0146: o_data_a = 16'b1110110000010000;
            14'h0147: o_data_a = 16'b0000000000001110;
            14'h0148: o_data_a = 16'b1110001100001000;
            14'h0149: o_data_a = 16'b0000000101001101;
            14'h014a: o_data_a = 16'b1110110000010000;
            14'h014b: o_data_a = 16'b0000000001011111;
            14'h014c: o_data_a = 16'b1110101010000111;
            14'h014d: o_data_a = 16'b0000000000000000;
            14'h014e: o_data_a = 16'b1111110010101000;
            14'h014f: o_data_a = 16'b1111110000010000;
            14'h0150: o_data_a = 16'b0000000000000101;
            14'h0151: o_data_a = 16'b1110001100001000;
            14'h0152: o_data_a = 16'b0000000000000011;
            14'h0153: o_data_a = 16'b1111110000010000;
            14'h0154: o_data_a = 16'b0000000000000000;
            14'h0155: o_data_a = 16'b1111110111101000;
            14'h0156: o_data_a = 16'b1110110010100000;
            14'h0157: o_data_a = 16'b1110001100001000;
            14'h0158: o_data_a = 16'b0000000000110110;
            14'h0159: o_data_a = 16'b1110101010000111;
            14'h015a: o_data_a = 16'b0000000000000010;
            14'h015b: o_data_a = 16'b1111110000100000;
            14'h015c: o_data_a = 16'b1111110000010000;
            14'h015d: o_data_a = 16'b0000000000000000;
            14'h015e: o_data_a = 16'b1111110111101000;
            14'h015f: o_data_a = 16'b1110110010100000;
            14'h0160: o_data_a = 16'b1110001100001000;
            14'h0161: o_data_a = 16'b0000000000000000;
            14'h0162: o_data_a = 16'b1111110010101000;
            14'h0163: o_data_a = 16'b1111110000010000;
            14'h0164: o_data_a = 16'b0000000000000011;
            14'h0165: o_data_a = 16'b1110001100001000;
            14'h0166: o_data_a = 16'b0000000000000011;
            14'h0167: o_data_a = 16'b1111110000010000;
            14'h0168: o_data_a = 16'b0000000000000000;
            14'h0169: o_data_a = 16'b1111110111101000;
            14'h016a: o_data_a = 16'b1110110010100000;
            14'h016b: o_data_a = 16'b1110001100001000;
            14'h016c: o_data_a = 16'b0000000000000001;
            14'h016d: o_data_a = 16'b1110110000010000;
            14'h016e: o_data_a = 16'b0000000000001101;
            14'h016f: o_data_a = 16'b1110001100001000;
            14'h0170: o_data_a = 16'b0010010010001101;
            14'h0171: o_data_a = 16'b1110110000010000;
            14'h0172: o_data_a = 16'b0000000000001110;
            14'h0173: o_data_a = 16'b1110001100001000;
            14'h0174: o_data_a = 16'b0000000101111000;
            14'h0175: o_data_a = 16'b1110110000010000;
            14'h0176: o_data_a = 16'b0000000001011111;
            14'h0177: o_data_a = 16'b1110101010000111;
            14'h0178: o_data_a = 16'b0000000000000000;
            14'h0179: o_data_a = 16'b1111110010101000;
            14'h017a: o_data_a = 16'b1111110000010000;
            14'h017b: o_data_a = 16'b0000000000000101;
            14'h017c: o_data_a = 16'b1110001100001000;
            14'h017d: o_data_a = 16'b0000000000000000;
            14'h017e: o_data_a = 16'b1111110111001000;
            14'h017f: o_data_a = 16'b1111110010100000;
            14'h0180: o_data_a = 16'b1110101010001000;
            14'h0181: o_data_a = 16'b0000000000110110;
            14'h0182: o_data_a = 16'b1110101010000111;
            14'h0183: o_data_a = 16'b0000000000000010;
            14'h0184: o_data_a = 16'b1111110000100000;
            14'h0185: o_data_a = 16'b1111110000010000;
            14'h0186: o_data_a = 16'b0000000000000000;
            14'h0187: o_data_a = 16'b1111110111101000;
            14'h0188: o_data_a = 16'b1110110010100000;
            14'h0189: o_data_a = 16'b1110001100001000;
            14'h018a: o_data_a = 16'b0000000000000000;
            14'h018b: o_data_a = 16'b1111110010101000;
            14'h018c: o_data_a = 16'b1111110000010000;
            14'h018d: o_data_a = 16'b0000000000000011;
            14'h018e: o_data_a = 16'b1110001100001000;
            14'h018f: o_data_a = 16'b0000000000000000;
            14'h0190: o_data_a = 16'b1111110111001000;
            14'h0191: o_data_a = 16'b1111110010100000;
            14'h0192: o_data_a = 16'b1110101010001000;
            14'h0193: o_data_a = 16'b0000000000000000;
            14'h0194: o_data_a = 16'b1111110010100000;
            14'h0195: o_data_a = 16'b1111110001001000;
            14'h0196: o_data_a = 16'b0000000000000001;
            14'h0197: o_data_a = 16'b1110110000010000;
            14'h0198: o_data_a = 16'b0000000000001101;
            14'h0199: o_data_a = 16'b1110001100001000;
            14'h019a: o_data_a = 16'b0101000110011001;
            14'h019b: o_data_a = 16'b1110110000010000;
            14'h019c: o_data_a = 16'b0000000000001110;
            14'h019d: o_data_a = 16'b1110001100001000;
            14'h019e: o_data_a = 16'b0000000110100010;
            14'h019f: o_data_a = 16'b1110110000010000;
            14'h01a0: o_data_a = 16'b0000000001011111;
            14'h01a1: o_data_a = 16'b1110101010000111;
            14'h01a2: o_data_a = 16'b0000000000000000;
            14'h01a3: o_data_a = 16'b1111110010101000;
            14'h01a4: o_data_a = 16'b1111110000010000;
            14'h01a5: o_data_a = 16'b0000000000000101;
            14'h01a6: o_data_a = 16'b1110001100001000;
            14'h01a7: o_data_a = 16'b0000000000000011;
            14'h01a8: o_data_a = 16'b1111110000010000;
            14'h01a9: o_data_a = 16'b0000000000000000;
            14'h01aa: o_data_a = 16'b1111110111101000;
            14'h01ab: o_data_a = 16'b1110110010100000;
            14'h01ac: o_data_a = 16'b1110001100001000;
            14'h01ad: o_data_a = 16'b0000000000000001;
            14'h01ae: o_data_a = 16'b1110110000010000;
            14'h01af: o_data_a = 16'b0000000000001101;
            14'h01b0: o_data_a = 16'b1110001100001000;
            14'h01b1: o_data_a = 16'b0000001000000010;
            14'h01b2: o_data_a = 16'b1110110000010000;
            14'h01b3: o_data_a = 16'b0000000000001110;
            14'h01b4: o_data_a = 16'b1110001100001000;
            14'h01b5: o_data_a = 16'b0000000110111001;
            14'h01b6: o_data_a = 16'b1110110000010000;
            14'h01b7: o_data_a = 16'b0000000001011111;
            14'h01b8: o_data_a = 16'b1110101010000111;
            14'h01b9: o_data_a = 16'b0000000000000000;
            14'h01ba: o_data_a = 16'b1111110010101000;
            14'h01bb: o_data_a = 16'b1111110000010000;
            14'h01bc: o_data_a = 16'b0000000000000101;
            14'h01bd: o_data_a = 16'b1110001100001000;
            14'h01be: o_data_a = 16'b0000000000000000;
            14'h01bf: o_data_a = 16'b1111110111001000;
            14'h01c0: o_data_a = 16'b1111110010100000;
            14'h01c1: o_data_a = 16'b1110101010001000;
            14'h01c2: o_data_a = 16'b0000000000110110;
            14'h01c3: o_data_a = 16'b1110101010000111;
            14'h01c4: o_data_a = 16'b0000000000000010;
            14'h01c5: o_data_a = 16'b1111110000100000;
            14'h01c6: o_data_a = 16'b1111110000010000;
            14'h01c7: o_data_a = 16'b0000000000000000;
            14'h01c8: o_data_a = 16'b1111110111101000;
            14'h01c9: o_data_a = 16'b1110110010100000;
            14'h01ca: o_data_a = 16'b1110001100001000;
            14'h01cb: o_data_a = 16'b0000000000000000;
            14'h01cc: o_data_a = 16'b1111110010101000;
            14'h01cd: o_data_a = 16'b1111110000010000;
            14'h01ce: o_data_a = 16'b0000000000000011;
            14'h01cf: o_data_a = 16'b1110001100001000;
            14'h01d0: o_data_a = 16'b0000000000000000;
            14'h01d1: o_data_a = 16'b1111110111001000;
            14'h01d2: o_data_a = 16'b1111110010100000;
            14'h01d3: o_data_a = 16'b1110101010001000;
            14'h01d4: o_data_a = 16'b0000000000000001;
            14'h01d5: o_data_a = 16'b1110110000010000;
            14'h01d6: o_data_a = 16'b0000000000001101;
            14'h01d7: o_data_a = 16'b1110001100001000;
            14'h01d8: o_data_a = 16'b0101000110011001;
            14'h01d9: o_data_a = 16'b1110110000010000;
            14'h01da: o_data_a = 16'b0000000000001110;
            14'h01db: o_data_a = 16'b1110001100001000;
            14'h01dc: o_data_a = 16'b0000000111100000;
            14'h01dd: o_data_a = 16'b1110110000010000;
            14'h01de: o_data_a = 16'b0000000001011111;
            14'h01df: o_data_a = 16'b1110101010000111;
            14'h01e0: o_data_a = 16'b0000000000000000;
            14'h01e1: o_data_a = 16'b1111110010101000;
            14'h01e2: o_data_a = 16'b1111110000010000;
            14'h01e3: o_data_a = 16'b0000000000000101;
            14'h01e4: o_data_a = 16'b1110001100001000;
            14'h01e5: o_data_a = 16'b0000000000000011;
            14'h01e6: o_data_a = 16'b1111110000010000;
            14'h01e7: o_data_a = 16'b0000000000000000;
            14'h01e8: o_data_a = 16'b1111110111101000;
            14'h01e9: o_data_a = 16'b1110110010100000;
            14'h01ea: o_data_a = 16'b1110001100001000;
            14'h01eb: o_data_a = 16'b0000000000000001;
            14'h01ec: o_data_a = 16'b1110110000010000;
            14'h01ed: o_data_a = 16'b0000000000001101;
            14'h01ee: o_data_a = 16'b1110001100001000;
            14'h01ef: o_data_a = 16'b0000001000000010;
            14'h01f0: o_data_a = 16'b1110110000010000;
            14'h01f1: o_data_a = 16'b0000000000001110;
            14'h01f2: o_data_a = 16'b1110001100001000;
            14'h01f3: o_data_a = 16'b0000000111110111;
            14'h01f4: o_data_a = 16'b1110110000010000;
            14'h01f5: o_data_a = 16'b0000000001011111;
            14'h01f6: o_data_a = 16'b1110101010000111;
            14'h01f7: o_data_a = 16'b0000000000000000;
            14'h01f8: o_data_a = 16'b1111110010101000;
            14'h01f9: o_data_a = 16'b1111110000010000;
            14'h01fa: o_data_a = 16'b0000000000000101;
            14'h01fb: o_data_a = 16'b1110001100001000;
            14'h01fc: o_data_a = 16'b0000000000000000;
            14'h01fd: o_data_a = 16'b1111110111001000;
            14'h01fe: o_data_a = 16'b1111110010100000;
            14'h01ff: o_data_a = 16'b1110101010001000;
            14'h0200: o_data_a = 16'b0000000000110110;
            14'h0201: o_data_a = 16'b1110101010000111;
            14'h0202: o_data_a = 16'b0000000000000010;
            14'h0203: o_data_a = 16'b1111110000100000;
            14'h0204: o_data_a = 16'b1111110000010000;
            14'h0205: o_data_a = 16'b0000000000000000;
            14'h0206: o_data_a = 16'b1111110111101000;
            14'h0207: o_data_a = 16'b1110110010100000;
            14'h0208: o_data_a = 16'b1110001100001000;
            14'h0209: o_data_a = 16'b0000000000000000;
            14'h020a: o_data_a = 16'b1111110010101000;
            14'h020b: o_data_a = 16'b1111110000010000;
            14'h020c: o_data_a = 16'b0000000000000011;
            14'h020d: o_data_a = 16'b1110001100001000;
            14'h020e: o_data_a = 16'b0000000000000011;
            14'h020f: o_data_a = 16'b1111110000100000;
            14'h0210: o_data_a = 16'b1111110000010000;
            14'h0211: o_data_a = 16'b0000000000000000;
            14'h0212: o_data_a = 16'b1111110111101000;
            14'h0213: o_data_a = 16'b1110110010100000;
            14'h0214: o_data_a = 16'b1110001100001000;
            14'h0215: o_data_a = 16'b0000000000000011;
            14'h0216: o_data_a = 16'b1111110111100000;
            14'h0217: o_data_a = 16'b1111110000010000;
            14'h0218: o_data_a = 16'b0000000000000000;
            14'h0219: o_data_a = 16'b1111110111101000;
            14'h021a: o_data_a = 16'b1110110010100000;
            14'h021b: o_data_a = 16'b1110001100001000;
            14'h021c: o_data_a = 16'b0000000000000011;
            14'h021d: o_data_a = 16'b1111110000100000;
            14'h021e: o_data_a = 16'b1111110000010000;
            14'h021f: o_data_a = 16'b0000000000000000;
            14'h0220: o_data_a = 16'b1111110111101000;
            14'h0221: o_data_a = 16'b1110110010100000;
            14'h0222: o_data_a = 16'b1110001100001000;
            14'h0223: o_data_a = 16'b0000000000000101;
            14'h0224: o_data_a = 16'b1110110000010000;
            14'h0225: o_data_a = 16'b0000000000000000;
            14'h0226: o_data_a = 16'b1111110111101000;
            14'h0227: o_data_a = 16'b1110110010100000;
            14'h0228: o_data_a = 16'b1110001100001000;
            14'h0229: o_data_a = 16'b0000000000000000;
            14'h022a: o_data_a = 16'b1111110010101000;
            14'h022b: o_data_a = 16'b1111110000010000;
            14'h022c: o_data_a = 16'b1110110010100000;
            14'h022d: o_data_a = 16'b1111000010001000;
            14'h022e: o_data_a = 16'b0000000000000011;
            14'h022f: o_data_a = 16'b1111110111100000;
            14'h0230: o_data_a = 16'b1111110000010000;
            14'h0231: o_data_a = 16'b0000000000000000;
            14'h0232: o_data_a = 16'b1111110111101000;
            14'h0233: o_data_a = 16'b1110110010100000;
            14'h0234: o_data_a = 16'b1110001100001000;
            14'h0235: o_data_a = 16'b0000000000000101;
            14'h0236: o_data_a = 16'b1110110000010000;
            14'h0237: o_data_a = 16'b0000000000000000;
            14'h0238: o_data_a = 16'b1111110111101000;
            14'h0239: o_data_a = 16'b1110110010100000;
            14'h023a: o_data_a = 16'b1110001100001000;
            14'h023b: o_data_a = 16'b0000000000000000;
            14'h023c: o_data_a = 16'b1111110010101000;
            14'h023d: o_data_a = 16'b1111110000010000;
            14'h023e: o_data_a = 16'b1110110010100000;
            14'h023f: o_data_a = 16'b1111000010001000;
            14'h0240: o_data_a = 16'b0000000000000100;
            14'h0241: o_data_a = 16'b1110110000010000;
            14'h0242: o_data_a = 16'b0000000000001101;
            14'h0243: o_data_a = 16'b1110001100001000;
            14'h0244: o_data_a = 16'b0101011101010010;
            14'h0245: o_data_a = 16'b1110110000010000;
            14'h0246: o_data_a = 16'b0000000000001110;
            14'h0247: o_data_a = 16'b1110001100001000;
            14'h0248: o_data_a = 16'b0000001001001100;
            14'h0249: o_data_a = 16'b1110110000010000;
            14'h024a: o_data_a = 16'b0000000001011111;
            14'h024b: o_data_a = 16'b1110101010000111;
            14'h024c: o_data_a = 16'b0000000000000000;
            14'h024d: o_data_a = 16'b1111110010101000;
            14'h024e: o_data_a = 16'b1111110000010000;
            14'h024f: o_data_a = 16'b0000000000000101;
            14'h0250: o_data_a = 16'b1110001100001000;
            14'h0251: o_data_a = 16'b0000000000000000;
            14'h0252: o_data_a = 16'b1111110111001000;
            14'h0253: o_data_a = 16'b1111110010100000;
            14'h0254: o_data_a = 16'b1110101010001000;
            14'h0255: o_data_a = 16'b0000000000110110;
            14'h0256: o_data_a = 16'b1110101010000111;
            14'h0257: o_data_a = 16'b0000000000000010;
            14'h0258: o_data_a = 16'b1111110000100000;
            14'h0259: o_data_a = 16'b1111110000010000;
            14'h025a: o_data_a = 16'b0000000000000000;
            14'h025b: o_data_a = 16'b1111110111101000;
            14'h025c: o_data_a = 16'b1110110010100000;
            14'h025d: o_data_a = 16'b1110001100001000;
            14'h025e: o_data_a = 16'b0000000000000000;
            14'h025f: o_data_a = 16'b1111110010101000;
            14'h0260: o_data_a = 16'b1111110000010000;
            14'h0261: o_data_a = 16'b0000000000000011;
            14'h0262: o_data_a = 16'b1110001100001000;
            14'h0263: o_data_a = 16'b0000000000000011;
            14'h0264: o_data_a = 16'b1111110000100000;
            14'h0265: o_data_a = 16'b1111110000010000;
            14'h0266: o_data_a = 16'b0000000000000000;
            14'h0267: o_data_a = 16'b1111110111101000;
            14'h0268: o_data_a = 16'b1110110010100000;
            14'h0269: o_data_a = 16'b1110001100001000;
            14'h026a: o_data_a = 16'b0000000000110110;
            14'h026b: o_data_a = 16'b1110101010000111;
            14'h026c: o_data_a = 16'b0000000000000010;
            14'h026d: o_data_a = 16'b1111110000100000;
            14'h026e: o_data_a = 16'b1111110000010000;
            14'h026f: o_data_a = 16'b0000000000000000;
            14'h0270: o_data_a = 16'b1111110111101000;
            14'h0271: o_data_a = 16'b1110110010100000;
            14'h0272: o_data_a = 16'b1110001100001000;
            14'h0273: o_data_a = 16'b0000000000000000;
            14'h0274: o_data_a = 16'b1111110010101000;
            14'h0275: o_data_a = 16'b1111110000010000;
            14'h0276: o_data_a = 16'b0000000000000011;
            14'h0277: o_data_a = 16'b1110001100001000;
            14'h0278: o_data_a = 16'b0000000000000011;
            14'h0279: o_data_a = 16'b1111110000100000;
            14'h027a: o_data_a = 16'b1111110000010000;
            14'h027b: o_data_a = 16'b0000000000000000;
            14'h027c: o_data_a = 16'b1111110111101000;
            14'h027d: o_data_a = 16'b1110110010100000;
            14'h027e: o_data_a = 16'b1110001100001000;
            14'h027f: o_data_a = 16'b0000000000000101;
            14'h0280: o_data_a = 16'b1110110000010000;
            14'h0281: o_data_a = 16'b0000000000000000;
            14'h0282: o_data_a = 16'b1111110111101000;
            14'h0283: o_data_a = 16'b1110110010100000;
            14'h0284: o_data_a = 16'b1110001100001000;
            14'h0285: o_data_a = 16'b0000000000000000;
            14'h0286: o_data_a = 16'b1111110010101000;
            14'h0287: o_data_a = 16'b1111110000010000;
            14'h0288: o_data_a = 16'b1110110010100000;
            14'h0289: o_data_a = 16'b1111000010001000;
            14'h028a: o_data_a = 16'b0000000000110110;
            14'h028b: o_data_a = 16'b1110101010000111;
            14'h028c: o_data_a = 16'b0000000000000011;
            14'h028d: o_data_a = 16'b1110110000010000;
            14'h028e: o_data_a = 16'b1110001110010000;
            14'h028f: o_data_a = 16'b0000000000000000;
            14'h0290: o_data_a = 16'b1111110111101000;
            14'h0291: o_data_a = 16'b1110110010100000;
            14'h0292: o_data_a = 16'b1110101010001000;
            14'h0293: o_data_a = 16'b0000001010001110;
            14'h0294: o_data_a = 16'b1110001100000001;
            14'h0295: o_data_a = 16'b0000000000000010;
            14'h0296: o_data_a = 16'b1111110000100000;
            14'h0297: o_data_a = 16'b1111110000010000;
            14'h0298: o_data_a = 16'b0000000000000000;
            14'h0299: o_data_a = 16'b1111110111101000;
            14'h029a: o_data_a = 16'b1110110010100000;
            14'h029b: o_data_a = 16'b1110001100001000;
            14'h029c: o_data_a = 16'b0000000000000000;
            14'h029d: o_data_a = 16'b1111110010101000;
            14'h029e: o_data_a = 16'b1111110000010000;
            14'h029f: o_data_a = 16'b0000000000000011;
            14'h02a0: o_data_a = 16'b1110001100001000;
            14'h02a1: o_data_a = 16'b0000000000000010;
            14'h02a2: o_data_a = 16'b1111110111100000;
            14'h02a3: o_data_a = 16'b1111110000010000;
            14'h02a4: o_data_a = 16'b0000000000000000;
            14'h02a5: o_data_a = 16'b1111110111101000;
            14'h02a6: o_data_a = 16'b1110110010100000;
            14'h02a7: o_data_a = 16'b1110001100001000;
            14'h02a8: o_data_a = 16'b0000000000000011;
            14'h02a9: o_data_a = 16'b1111110000100000;
            14'h02aa: o_data_a = 16'b1111110000010000;
            14'h02ab: o_data_a = 16'b0000000000000000;
            14'h02ac: o_data_a = 16'b1111110111101000;
            14'h02ad: o_data_a = 16'b1110110010100000;
            14'h02ae: o_data_a = 16'b1110001100001000;
            14'h02af: o_data_a = 16'b0000000000000000;
            14'h02b0: o_data_a = 16'b1111110010101000;
            14'h02b1: o_data_a = 16'b1111110000010000;
            14'h02b2: o_data_a = 16'b1110110010100000;
            14'h02b3: o_data_a = 16'b1111000111001000;
            14'h02b4: o_data_a = 16'b0000000000000000;
            14'h02b5: o_data_a = 16'b1111110010101000;
            14'h02b6: o_data_a = 16'b1111110000010000;
            14'h02b7: o_data_a = 16'b0000000000000011;
            14'h02b8: o_data_a = 16'b1111110111100000;
            14'h02b9: o_data_a = 16'b1110110111100000;
            14'h02ba: o_data_a = 16'b1110001100001000;
            14'h02bb: o_data_a = 16'b0000000000000010;
            14'h02bc: o_data_a = 16'b1111110111100000;
            14'h02bd: o_data_a = 16'b1110110111100000;
            14'h02be: o_data_a = 16'b1111110000010000;
            14'h02bf: o_data_a = 16'b0000000000000000;
            14'h02c0: o_data_a = 16'b1111110111101000;
            14'h02c1: o_data_a = 16'b1110110010100000;
            14'h02c2: o_data_a = 16'b1110001100001000;
            14'h02c3: o_data_a = 16'b0000000000000011;
            14'h02c4: o_data_a = 16'b1111110111100000;
            14'h02c5: o_data_a = 16'b1111110000010000;
            14'h02c6: o_data_a = 16'b0000000000000000;
            14'h02c7: o_data_a = 16'b1111110111101000;
            14'h02c8: o_data_a = 16'b1110110010100000;
            14'h02c9: o_data_a = 16'b1110001100001000;
            14'h02ca: o_data_a = 16'b0000000000000000;
            14'h02cb: o_data_a = 16'b1111110010101000;
            14'h02cc: o_data_a = 16'b1111110000010000;
            14'h02cd: o_data_a = 16'b1110110010100000;
            14'h02ce: o_data_a = 16'b1111000111001000;
            14'h02cf: o_data_a = 16'b0000000000000000;
            14'h02d0: o_data_a = 16'b1111110010101000;
            14'h02d1: o_data_a = 16'b1111110000010000;
            14'h02d2: o_data_a = 16'b0000000000000011;
            14'h02d3: o_data_a = 16'b1111110111100000;
            14'h02d4: o_data_a = 16'b1110110111100000;
            14'h02d5: o_data_a = 16'b1110110111100000;
            14'h02d6: o_data_a = 16'b1110001100001000;
            14'h02d7: o_data_a = 16'b0000000000000011;
            14'h02d8: o_data_a = 16'b1111110111100000;
            14'h02d9: o_data_a = 16'b1110110111100000;
            14'h02da: o_data_a = 16'b1111110000010000;
            14'h02db: o_data_a = 16'b0000000000000000;
            14'h02dc: o_data_a = 16'b1111110111101000;
            14'h02dd: o_data_a = 16'b1110110010100000;
            14'h02de: o_data_a = 16'b1110001100001000;
            14'h02df: o_data_a = 16'b0000000000000001;
            14'h02e0: o_data_a = 16'b1110110000010000;
            14'h02e1: o_data_a = 16'b0000000000001101;
            14'h02e2: o_data_a = 16'b1110001100001000;
            14'h02e3: o_data_a = 16'b0001101001110110;
            14'h02e4: o_data_a = 16'b1110110000010000;
            14'h02e5: o_data_a = 16'b0000000000001110;
            14'h02e6: o_data_a = 16'b1110001100001000;
            14'h02e7: o_data_a = 16'b0000001011101011;
            14'h02e8: o_data_a = 16'b1110110000010000;
            14'h02e9: o_data_a = 16'b0000000001011111;
            14'h02ea: o_data_a = 16'b1110101010000111;
            14'h02eb: o_data_a = 16'b0000000000000000;
            14'h02ec: o_data_a = 16'b1111110010101000;
            14'h02ed: o_data_a = 16'b1111110000010000;
            14'h02ee: o_data_a = 16'b0000000000000001;
            14'h02ef: o_data_a = 16'b1111110000100000;
            14'h02f0: o_data_a = 16'b1110001100001000;
            14'h02f1: o_data_a = 16'b0000000000000011;
            14'h02f2: o_data_a = 16'b1111110000010000;
            14'h02f3: o_data_a = 16'b0000000000000011;
            14'h02f4: o_data_a = 16'b1110000010100000;
            14'h02f5: o_data_a = 16'b1111110000010000;
            14'h02f6: o_data_a = 16'b0000000000000000;
            14'h02f7: o_data_a = 16'b1111110111101000;
            14'h02f8: o_data_a = 16'b1110110010100000;
            14'h02f9: o_data_a = 16'b1110001100001000;
            14'h02fa: o_data_a = 16'b0000000000000001;
            14'h02fb: o_data_a = 16'b1110110000010000;
            14'h02fc: o_data_a = 16'b0000000000001101;
            14'h02fd: o_data_a = 16'b1110001100001000;
            14'h02fe: o_data_a = 16'b0001101001110110;
            14'h02ff: o_data_a = 16'b1110110000010000;
            14'h0300: o_data_a = 16'b0000000000001110;
            14'h0301: o_data_a = 16'b1110001100001000;
            14'h0302: o_data_a = 16'b0000001100000110;
            14'h0303: o_data_a = 16'b1110110000010000;
            14'h0304: o_data_a = 16'b0000000001011111;
            14'h0305: o_data_a = 16'b1110101010000111;
            14'h0306: o_data_a = 16'b0000000000000000;
            14'h0307: o_data_a = 16'b1111110010101000;
            14'h0308: o_data_a = 16'b1111110000010000;
            14'h0309: o_data_a = 16'b0000000000000001;
            14'h030a: o_data_a = 16'b1111110111100000;
            14'h030b: o_data_a = 16'b1110001100001000;
            14'h030c: o_data_a = 16'b0000000000000001;
            14'h030d: o_data_a = 16'b1111110000100000;
            14'h030e: o_data_a = 16'b1111110000010000;
            14'h030f: o_data_a = 16'b0000000000000000;
            14'h0310: o_data_a = 16'b1111110111101000;
            14'h0311: o_data_a = 16'b1110110010100000;
            14'h0312: o_data_a = 16'b1110001100001000;
            14'h0313: o_data_a = 16'b0000000000000001;
            14'h0314: o_data_a = 16'b1111110111100000;
            14'h0315: o_data_a = 16'b1111110000010000;
            14'h0316: o_data_a = 16'b0000000000000000;
            14'h0317: o_data_a = 16'b1111110111101000;
            14'h0318: o_data_a = 16'b1110110010100000;
            14'h0319: o_data_a = 16'b1110001100001000;
            14'h031a: o_data_a = 16'b0000001100011110;
            14'h031b: o_data_a = 16'b1110110000010000;
            14'h031c: o_data_a = 16'b0000000000100110;
            14'h031d: o_data_a = 16'b1110101010000111;
            14'h031e: o_data_a = 16'b0000000000000011;
            14'h031f: o_data_a = 16'b1111110000010000;
            14'h0320: o_data_a = 16'b0000000000000111;
            14'h0321: o_data_a = 16'b1110000010010000;
            14'h0322: o_data_a = 16'b0000000000001101;
            14'h0323: o_data_a = 16'b1110001100001000;
            14'h0324: o_data_a = 16'b0000000000000000;
            14'h0325: o_data_a = 16'b1111110010101000;
            14'h0326: o_data_a = 16'b1111110000010000;
            14'h0327: o_data_a = 16'b0000000000001101;
            14'h0328: o_data_a = 16'b1111110000100000;
            14'h0329: o_data_a = 16'b1110001100001000;
            14'h032a: o_data_a = 16'b0000000000000011;
            14'h032b: o_data_a = 16'b1111110000010000;
            14'h032c: o_data_a = 16'b0000000000000111;
            14'h032d: o_data_a = 16'b1110000010100000;
            14'h032e: o_data_a = 16'b1111110000010000;
            14'h032f: o_data_a = 16'b0000000000000000;
            14'h0330: o_data_a = 16'b1111110111101000;
            14'h0331: o_data_a = 16'b1110110010100000;
            14'h0332: o_data_a = 16'b1110001100001000;
            14'h0333: o_data_a = 16'b0000000000000000;
            14'h0334: o_data_a = 16'b1111110010101000;
            14'h0335: o_data_a = 16'b1111110000010000;
            14'h0336: o_data_a = 16'b0000001100111010;
            14'h0337: o_data_a = 16'b1110001100000101;
            14'h0338: o_data_a = 16'b0000001110100010;
            14'h0339: o_data_a = 16'b1110101010000111;
            14'h033a: o_data_a = 16'b0000000000000001;
            14'h033b: o_data_a = 16'b1111110000100000;
            14'h033c: o_data_a = 16'b1111110000010000;
            14'h033d: o_data_a = 16'b0000000000000000;
            14'h033e: o_data_a = 16'b1111110111101000;
            14'h033f: o_data_a = 16'b1110110010100000;
            14'h0340: o_data_a = 16'b1110001100001000;
            14'h0341: o_data_a = 16'b0000000000000000;
            14'h0342: o_data_a = 16'b1111110010101000;
            14'h0343: o_data_a = 16'b1111110000010000;
            14'h0344: o_data_a = 16'b0000000000000001;
            14'h0345: o_data_a = 16'b1111110111100000;
            14'h0346: o_data_a = 16'b1110110111100000;
            14'h0347: o_data_a = 16'b1110001100001000;
            14'h0348: o_data_a = 16'b0000000000000001;
            14'h0349: o_data_a = 16'b1111110111100000;
            14'h034a: o_data_a = 16'b1111110000010000;
            14'h034b: o_data_a = 16'b0000000000000000;
            14'h034c: o_data_a = 16'b1111110111101000;
            14'h034d: o_data_a = 16'b1110110010100000;
            14'h034e: o_data_a = 16'b1110001100001000;
            14'h034f: o_data_a = 16'b0000000000000000;
            14'h0350: o_data_a = 16'b1111110010101000;
            14'h0351: o_data_a = 16'b1111110000010000;
            14'h0352: o_data_a = 16'b0000000000000001;
            14'h0353: o_data_a = 16'b1111110000100000;
            14'h0354: o_data_a = 16'b1110001100001000;
            14'h0355: o_data_a = 16'b0000000000000001;
            14'h0356: o_data_a = 16'b1111110111100000;
            14'h0357: o_data_a = 16'b1110110111100000;
            14'h0358: o_data_a = 16'b1111110000010000;
            14'h0359: o_data_a = 16'b0000000000000000;
            14'h035a: o_data_a = 16'b1111110111101000;
            14'h035b: o_data_a = 16'b1110110010100000;
            14'h035c: o_data_a = 16'b1110001100001000;
            14'h035d: o_data_a = 16'b0000000000000000;
            14'h035e: o_data_a = 16'b1111110010101000;
            14'h035f: o_data_a = 16'b1111110000010000;
            14'h0360: o_data_a = 16'b0000000000000001;
            14'h0361: o_data_a = 16'b1111110111100000;
            14'h0362: o_data_a = 16'b1110001100001000;
            14'h0363: o_data_a = 16'b0000000000000011;
            14'h0364: o_data_a = 16'b1111110111100000;
            14'h0365: o_data_a = 16'b1111110000010000;
            14'h0366: o_data_a = 16'b0000000000000000;
            14'h0367: o_data_a = 16'b1111110111101000;
            14'h0368: o_data_a = 16'b1110110010100000;
            14'h0369: o_data_a = 16'b1110001100001000;
            14'h036a: o_data_a = 16'b0000000000000010;
            14'h036b: o_data_a = 16'b1111110111100000;
            14'h036c: o_data_a = 16'b1110110111100000;
            14'h036d: o_data_a = 16'b1111110000010000;
            14'h036e: o_data_a = 16'b0000000000000000;
            14'h036f: o_data_a = 16'b1111110111101000;
            14'h0370: o_data_a = 16'b1110110010100000;
            14'h0371: o_data_a = 16'b1110001100001000;
            14'h0372: o_data_a = 16'b0000001101110110;
            14'h0373: o_data_a = 16'b1110110000010000;
            14'h0374: o_data_a = 16'b0000000000100110;
            14'h0375: o_data_a = 16'b1110101010000111;
            14'h0376: o_data_a = 16'b0000000000000011;
            14'h0377: o_data_a = 16'b1111110000010000;
            14'h0378: o_data_a = 16'b0000000000001000;
            14'h0379: o_data_a = 16'b1110000010010000;
            14'h037a: o_data_a = 16'b0000000000001101;
            14'h037b: o_data_a = 16'b1110001100001000;
            14'h037c: o_data_a = 16'b0000000000000000;
            14'h037d: o_data_a = 16'b1111110010101000;
            14'h037e: o_data_a = 16'b1111110000010000;
            14'h037f: o_data_a = 16'b0000000000001101;
            14'h0380: o_data_a = 16'b1111110000100000;
            14'h0381: o_data_a = 16'b1110001100001000;
            14'h0382: o_data_a = 16'b0000000000000011;
            14'h0383: o_data_a = 16'b1111110000100000;
            14'h0384: o_data_a = 16'b1111110000010000;
            14'h0385: o_data_a = 16'b0000000000000000;
            14'h0386: o_data_a = 16'b1111110111101000;
            14'h0387: o_data_a = 16'b1110110010100000;
            14'h0388: o_data_a = 16'b1110001100001000;
            14'h0389: o_data_a = 16'b0000000000000010;
            14'h038a: o_data_a = 16'b1111110111100000;
            14'h038b: o_data_a = 16'b1111110000010000;
            14'h038c: o_data_a = 16'b0000000000000000;
            14'h038d: o_data_a = 16'b1111110111101000;
            14'h038e: o_data_a = 16'b1110110010100000;
            14'h038f: o_data_a = 16'b1110001100001000;
            14'h0390: o_data_a = 16'b0000001110010100;
            14'h0391: o_data_a = 16'b1110110000010000;
            14'h0392: o_data_a = 16'b0000000000100110;
            14'h0393: o_data_a = 16'b1110101010000111;
            14'h0394: o_data_a = 16'b0000000000000011;
            14'h0395: o_data_a = 16'b1111110000010000;
            14'h0396: o_data_a = 16'b0000000000001001;
            14'h0397: o_data_a = 16'b1110000010010000;
            14'h0398: o_data_a = 16'b0000000000001101;
            14'h0399: o_data_a = 16'b1110001100001000;
            14'h039a: o_data_a = 16'b0000000000000000;
            14'h039b: o_data_a = 16'b1111110010101000;
            14'h039c: o_data_a = 16'b1111110000010000;
            14'h039d: o_data_a = 16'b0000000000001101;
            14'h039e: o_data_a = 16'b1111110000100000;
            14'h039f: o_data_a = 16'b1110001100001000;
            14'h03a0: o_data_a = 16'b0000001111011111;
            14'h03a1: o_data_a = 16'b1110101010000111;
            14'h03a2: o_data_a = 16'b0000000000000011;
            14'h03a3: o_data_a = 16'b1111110000100000;
            14'h03a4: o_data_a = 16'b1111110000010000;
            14'h03a5: o_data_a = 16'b0000000000000000;
            14'h03a6: o_data_a = 16'b1111110111101000;
            14'h03a7: o_data_a = 16'b1110110010100000;
            14'h03a8: o_data_a = 16'b1110001100001000;
            14'h03a9: o_data_a = 16'b0000000000000010;
            14'h03aa: o_data_a = 16'b1111110111100000;
            14'h03ab: o_data_a = 16'b1111110000010000;
            14'h03ac: o_data_a = 16'b0000000000000000;
            14'h03ad: o_data_a = 16'b1111110111101000;
            14'h03ae: o_data_a = 16'b1110110010100000;
            14'h03af: o_data_a = 16'b1110001100001000;
            14'h03b0: o_data_a = 16'b0000001110110100;
            14'h03b1: o_data_a = 16'b1110110000010000;
            14'h03b2: o_data_a = 16'b0000000000100110;
            14'h03b3: o_data_a = 16'b1110101010000111;
            14'h03b4: o_data_a = 16'b0000000000000011;
            14'h03b5: o_data_a = 16'b1111110000010000;
            14'h03b6: o_data_a = 16'b0000000000001000;
            14'h03b7: o_data_a = 16'b1110000010010000;
            14'h03b8: o_data_a = 16'b0000000000001101;
            14'h03b9: o_data_a = 16'b1110001100001000;
            14'h03ba: o_data_a = 16'b0000000000000000;
            14'h03bb: o_data_a = 16'b1111110010101000;
            14'h03bc: o_data_a = 16'b1111110000010000;
            14'h03bd: o_data_a = 16'b0000000000001101;
            14'h03be: o_data_a = 16'b1111110000100000;
            14'h03bf: o_data_a = 16'b1110001100001000;
            14'h03c0: o_data_a = 16'b0000000000000011;
            14'h03c1: o_data_a = 16'b1111110111100000;
            14'h03c2: o_data_a = 16'b1111110000010000;
            14'h03c3: o_data_a = 16'b0000000000000000;
            14'h03c4: o_data_a = 16'b1111110111101000;
            14'h03c5: o_data_a = 16'b1110110010100000;
            14'h03c6: o_data_a = 16'b1110001100001000;
            14'h03c7: o_data_a = 16'b0000000000000010;
            14'h03c8: o_data_a = 16'b1111110111100000;
            14'h03c9: o_data_a = 16'b1110110111100000;
            14'h03ca: o_data_a = 16'b1111110000010000;
            14'h03cb: o_data_a = 16'b0000000000000000;
            14'h03cc: o_data_a = 16'b1111110111101000;
            14'h03cd: o_data_a = 16'b1110110010100000;
            14'h03ce: o_data_a = 16'b1110001100001000;
            14'h03cf: o_data_a = 16'b0000001111010011;
            14'h03d0: o_data_a = 16'b1110110000010000;
            14'h03d1: o_data_a = 16'b0000000000100110;
            14'h03d2: o_data_a = 16'b1110101010000111;
            14'h03d3: o_data_a = 16'b0000000000000011;
            14'h03d4: o_data_a = 16'b1111110000010000;
            14'h03d5: o_data_a = 16'b0000000000001001;
            14'h03d6: o_data_a = 16'b1110000010010000;
            14'h03d7: o_data_a = 16'b0000000000001101;
            14'h03d8: o_data_a = 16'b1110001100001000;
            14'h03d9: o_data_a = 16'b0000000000000000;
            14'h03da: o_data_a = 16'b1111110010101000;
            14'h03db: o_data_a = 16'b1111110000010000;
            14'h03dc: o_data_a = 16'b0000000000001101;
            14'h03dd: o_data_a = 16'b1111110000100000;
            14'h03de: o_data_a = 16'b1110001100001000;
            14'h03df: o_data_a = 16'b0000000000000010;
            14'h03e0: o_data_a = 16'b1110110000010000;
            14'h03e1: o_data_a = 16'b0000000000000000;
            14'h03e2: o_data_a = 16'b1111110111101000;
            14'h03e3: o_data_a = 16'b1110110010100000;
            14'h03e4: o_data_a = 16'b1110001100001000;
            14'h03e5: o_data_a = 16'b0000000000000001;
            14'h03e6: o_data_a = 16'b1111110111100000;
            14'h03e7: o_data_a = 16'b1111110000010000;
            14'h03e8: o_data_a = 16'b0000000000000000;
            14'h03e9: o_data_a = 16'b1111110111101000;
            14'h03ea: o_data_a = 16'b1110110010100000;
            14'h03eb: o_data_a = 16'b1110001100001000;
            14'h03ec: o_data_a = 16'b0000000000000010;
            14'h03ed: o_data_a = 16'b1110110000010000;
            14'h03ee: o_data_a = 16'b0000000000001101;
            14'h03ef: o_data_a = 16'b1110001100001000;
            14'h03f0: o_data_a = 16'b0001101010100110;
            14'h03f1: o_data_a = 16'b1110110000010000;
            14'h03f2: o_data_a = 16'b0000000000001110;
            14'h03f3: o_data_a = 16'b1110001100001000;
            14'h03f4: o_data_a = 16'b0000001111111000;
            14'h03f5: o_data_a = 16'b1110110000010000;
            14'h03f6: o_data_a = 16'b0000000001011111;
            14'h03f7: o_data_a = 16'b1110101010000111;
            14'h03f8: o_data_a = 16'b0000000000000001;
            14'h03f9: o_data_a = 16'b1111110000100000;
            14'h03fa: o_data_a = 16'b1111110000010000;
            14'h03fb: o_data_a = 16'b0000000000000000;
            14'h03fc: o_data_a = 16'b1111110111101000;
            14'h03fd: o_data_a = 16'b1110110010100000;
            14'h03fe: o_data_a = 16'b1110001100001000;
            14'h03ff: o_data_a = 16'b0000000000000000;
            14'h0400: o_data_a = 16'b1111110010101000;
            14'h0401: o_data_a = 16'b1111110000010000;
            14'h0402: o_data_a = 16'b1110110010100000;
            14'h0403: o_data_a = 16'b1111000111001000;
            14'h0404: o_data_a = 16'b0000000000000000;
            14'h0405: o_data_a = 16'b1111110010101000;
            14'h0406: o_data_a = 16'b1111110000010000;
            14'h0407: o_data_a = 16'b0000000000000011;
            14'h0408: o_data_a = 16'b1111110111100000;
            14'h0409: o_data_a = 16'b1110110111100000;
            14'h040a: o_data_a = 16'b1110110111100000;
            14'h040b: o_data_a = 16'b1110110111100000;
            14'h040c: o_data_a = 16'b1110001100001000;
            14'h040d: o_data_a = 16'b0000000000000010;
            14'h040e: o_data_a = 16'b1110110000010000;
            14'h040f: o_data_a = 16'b0000000000000000;
            14'h0410: o_data_a = 16'b1111110111101000;
            14'h0411: o_data_a = 16'b1110110010100000;
            14'h0412: o_data_a = 16'b1110001100001000;
            14'h0413: o_data_a = 16'b0000000000000001;
            14'h0414: o_data_a = 16'b1111110111100000;
            14'h0415: o_data_a = 16'b1111110000010000;
            14'h0416: o_data_a = 16'b0000000000000000;
            14'h0417: o_data_a = 16'b1111110111101000;
            14'h0418: o_data_a = 16'b1110110010100000;
            14'h0419: o_data_a = 16'b1110001100001000;
            14'h041a: o_data_a = 16'b0000000000000010;
            14'h041b: o_data_a = 16'b1110110000010000;
            14'h041c: o_data_a = 16'b0000000000001101;
            14'h041d: o_data_a = 16'b1110001100001000;
            14'h041e: o_data_a = 16'b0001101010100110;
            14'h041f: o_data_a = 16'b1110110000010000;
            14'h0420: o_data_a = 16'b0000000000001110;
            14'h0421: o_data_a = 16'b1110001100001000;
            14'h0422: o_data_a = 16'b0000010000100110;
            14'h0423: o_data_a = 16'b1110110000010000;
            14'h0424: o_data_a = 16'b0000000001011111;
            14'h0425: o_data_a = 16'b1110101010000111;
            14'h0426: o_data_a = 16'b0000000000000000;
            14'h0427: o_data_a = 16'b1111110010101000;
            14'h0428: o_data_a = 16'b1111110000010000;
            14'h0429: o_data_a = 16'b0000000000000011;
            14'h042a: o_data_a = 16'b1111110111100000;
            14'h042b: o_data_a = 16'b1110110111100000;
            14'h042c: o_data_a = 16'b1110110111100000;
            14'h042d: o_data_a = 16'b1110110111100000;
            14'h042e: o_data_a = 16'b1110110111100000;
            14'h042f: o_data_a = 16'b1110001100001000;
            14'h0430: o_data_a = 16'b0000000000000010;
            14'h0431: o_data_a = 16'b1110110000010000;
            14'h0432: o_data_a = 16'b0000000000000000;
            14'h0433: o_data_a = 16'b1111110111101000;
            14'h0434: o_data_a = 16'b1110110010100000;
            14'h0435: o_data_a = 16'b1110001100001000;
            14'h0436: o_data_a = 16'b0000000000000001;
            14'h0437: o_data_a = 16'b1111110111100000;
            14'h0438: o_data_a = 16'b1111110000010000;
            14'h0439: o_data_a = 16'b0000000000000000;
            14'h043a: o_data_a = 16'b1111110111101000;
            14'h043b: o_data_a = 16'b1110110010100000;
            14'h043c: o_data_a = 16'b1110001100001000;
            14'h043d: o_data_a = 16'b0000000000000001;
            14'h043e: o_data_a = 16'b1111110000100000;
            14'h043f: o_data_a = 16'b1111110000010000;
            14'h0440: o_data_a = 16'b0000000000000000;
            14'h0441: o_data_a = 16'b1111110111101000;
            14'h0442: o_data_a = 16'b1110110010100000;
            14'h0443: o_data_a = 16'b1110001100001000;
            14'h0444: o_data_a = 16'b0000000000000000;
            14'h0445: o_data_a = 16'b1111110010101000;
            14'h0446: o_data_a = 16'b1111110000010000;
            14'h0447: o_data_a = 16'b1110110010100000;
            14'h0448: o_data_a = 16'b1111000111001000;
            14'h0449: o_data_a = 16'b0000000000000010;
            14'h044a: o_data_a = 16'b1110110000010000;
            14'h044b: o_data_a = 16'b0000000000001101;
            14'h044c: o_data_a = 16'b1110001100001000;
            14'h044d: o_data_a = 16'b0001101010100110;
            14'h044e: o_data_a = 16'b1110110000010000;
            14'h044f: o_data_a = 16'b0000000000001110;
            14'h0450: o_data_a = 16'b1110001100001000;
            14'h0451: o_data_a = 16'b0000010001010101;
            14'h0452: o_data_a = 16'b1110110000010000;
            14'h0453: o_data_a = 16'b0000000001011111;
            14'h0454: o_data_a = 16'b1110101010000111;
            14'h0455: o_data_a = 16'b0000000000000000;
            14'h0456: o_data_a = 16'b1111110010101000;
            14'h0457: o_data_a = 16'b1111110000010000;
            14'h0458: o_data_a = 16'b0000000000000011;
            14'h0459: o_data_a = 16'b1111110111100000;
            14'h045a: o_data_a = 16'b1110110111100000;
            14'h045b: o_data_a = 16'b1110110111100000;
            14'h045c: o_data_a = 16'b1110110111100000;
            14'h045d: o_data_a = 16'b1110110111100000;
            14'h045e: o_data_a = 16'b1110110111100000;
            14'h045f: o_data_a = 16'b1110001100001000;
            14'h0460: o_data_a = 16'b0000000000000000;
            14'h0461: o_data_a = 16'b1111110111001000;
            14'h0462: o_data_a = 16'b1111110010100000;
            14'h0463: o_data_a = 16'b1110101010001000;
            14'h0464: o_data_a = 16'b0000000000110110;
            14'h0465: o_data_a = 16'b1110101010000111;
            14'h0466: o_data_a = 16'b0000000000000010;
            14'h0467: o_data_a = 16'b1111110000100000;
            14'h0468: o_data_a = 16'b1111110000010000;
            14'h0469: o_data_a = 16'b0000000000000000;
            14'h046a: o_data_a = 16'b1111110111101000;
            14'h046b: o_data_a = 16'b1110110010100000;
            14'h046c: o_data_a = 16'b1110001100001000;
            14'h046d: o_data_a = 16'b0000000000000000;
            14'h046e: o_data_a = 16'b1111110010101000;
            14'h046f: o_data_a = 16'b1111110000010000;
            14'h0470: o_data_a = 16'b0000000000000011;
            14'h0471: o_data_a = 16'b1110001100001000;
            14'h0472: o_data_a = 16'b0000000000000011;
            14'h0473: o_data_a = 16'b1111110000010000;
            14'h0474: o_data_a = 16'b0000000000000000;
            14'h0475: o_data_a = 16'b1111110111101000;
            14'h0476: o_data_a = 16'b1110110010100000;
            14'h0477: o_data_a = 16'b1110001100001000;
            14'h0478: o_data_a = 16'b0000000000000001;
            14'h0479: o_data_a = 16'b1110110000010000;
            14'h047a: o_data_a = 16'b0000000000001101;
            14'h047b: o_data_a = 16'b1110001100001000;
            14'h047c: o_data_a = 16'b0000000111000100;
            14'h047d: o_data_a = 16'b1110110000010000;
            14'h047e: o_data_a = 16'b0000000000001110;
            14'h047f: o_data_a = 16'b1110001100001000;
            14'h0480: o_data_a = 16'b0000010010000100;
            14'h0481: o_data_a = 16'b1110110000010000;
            14'h0482: o_data_a = 16'b0000000001011111;
            14'h0483: o_data_a = 16'b1110101010000111;
            14'h0484: o_data_a = 16'b0000000000000000;
            14'h0485: o_data_a = 16'b1111110010101000;
            14'h0486: o_data_a = 16'b1111110000010000;
            14'h0487: o_data_a = 16'b0000000000000101;
            14'h0488: o_data_a = 16'b1110001100001000;
            14'h0489: o_data_a = 16'b0000000000000011;
            14'h048a: o_data_a = 16'b1111110000010000;
            14'h048b: o_data_a = 16'b0000000000000100;
            14'h048c: o_data_a = 16'b1110000010100000;
            14'h048d: o_data_a = 16'b1111110000010000;
            14'h048e: o_data_a = 16'b0000000000000000;
            14'h048f: o_data_a = 16'b1111110111101000;
            14'h0490: o_data_a = 16'b1110110010100000;
            14'h0491: o_data_a = 16'b1110001100001000;
            14'h0492: o_data_a = 16'b0000000000000000;
            14'h0493: o_data_a = 16'b1111110111001000;
            14'h0494: o_data_a = 16'b1111110010100000;
            14'h0495: o_data_a = 16'b1110101010001000;
            14'h0496: o_data_a = 16'b0000010010011010;
            14'h0497: o_data_a = 16'b1110110000010000;
            14'h0498: o_data_a = 16'b0000000000100110;
            14'h0499: o_data_a = 16'b1110101010000111;
            14'h049a: o_data_a = 16'b0000000000000000;
            14'h049b: o_data_a = 16'b1111110010101000;
            14'h049c: o_data_a = 16'b1111110000010000;
            14'h049d: o_data_a = 16'b0000010010100001;
            14'h049e: o_data_a = 16'b1110001100000101;
            14'h049f: o_data_a = 16'b0000010011000011;
            14'h04a0: o_data_a = 16'b1110101010000111;
            14'h04a1: o_data_a = 16'b0000000000000011;
            14'h04a2: o_data_a = 16'b1111110000010000;
            14'h04a3: o_data_a = 16'b0000000000000100;
            14'h04a4: o_data_a = 16'b1110000010100000;
            14'h04a5: o_data_a = 16'b1111110000010000;
            14'h04a6: o_data_a = 16'b0000000000000000;
            14'h04a7: o_data_a = 16'b1111110111101000;
            14'h04a8: o_data_a = 16'b1110110010100000;
            14'h04a9: o_data_a = 16'b1110001100001000;
            14'h04aa: o_data_a = 16'b0000000000000011;
            14'h04ab: o_data_a = 16'b1111110000010000;
            14'h04ac: o_data_a = 16'b0000000000000101;
            14'h04ad: o_data_a = 16'b1110000010100000;
            14'h04ae: o_data_a = 16'b1111110000010000;
            14'h04af: o_data_a = 16'b0000000000000000;
            14'h04b0: o_data_a = 16'b1111110111101000;
            14'h04b1: o_data_a = 16'b1110110010100000;
            14'h04b2: o_data_a = 16'b1110001100001000;
            14'h04b3: o_data_a = 16'b0000000000000000;
            14'h04b4: o_data_a = 16'b1111110010101000;
            14'h04b5: o_data_a = 16'b1111110000010000;
            14'h04b6: o_data_a = 16'b1110110010100000;
            14'h04b7: o_data_a = 16'b1111000010001000;
            14'h04b8: o_data_a = 16'b0000000000000000;
            14'h04b9: o_data_a = 16'b1111110010101000;
            14'h04ba: o_data_a = 16'b1111110000010000;
            14'h04bb: o_data_a = 16'b0000000000000011;
            14'h04bc: o_data_a = 16'b1111110111100000;
            14'h04bd: o_data_a = 16'b1110110111100000;
            14'h04be: o_data_a = 16'b1110110111100000;
            14'h04bf: o_data_a = 16'b1110110111100000;
            14'h04c0: o_data_a = 16'b1110001100001000;
            14'h04c1: o_data_a = 16'b0000010101111001;
            14'h04c2: o_data_a = 16'b1110101010000111;
            14'h04c3: o_data_a = 16'b0000000000000011;
            14'h04c4: o_data_a = 16'b1111110000010000;
            14'h04c5: o_data_a = 16'b0000000000000100;
            14'h04c6: o_data_a = 16'b1110000010100000;
            14'h04c7: o_data_a = 16'b1111110000010000;
            14'h04c8: o_data_a = 16'b0000000000000000;
            14'h04c9: o_data_a = 16'b1111110111101000;
            14'h04ca: o_data_a = 16'b1110110010100000;
            14'h04cb: o_data_a = 16'b1110001100001000;
            14'h04cc: o_data_a = 16'b0000000000000011;
            14'h04cd: o_data_a = 16'b1111110000010000;
            14'h04ce: o_data_a = 16'b0000000000000110;
            14'h04cf: o_data_a = 16'b1110000010100000;
            14'h04d0: o_data_a = 16'b1111110000010000;
            14'h04d1: o_data_a = 16'b0000000000000000;
            14'h04d2: o_data_a = 16'b1111110111101000;
            14'h04d3: o_data_a = 16'b1110110010100000;
            14'h04d4: o_data_a = 16'b1110001100001000;
            14'h04d5: o_data_a = 16'b0000000000000000;
            14'h04d6: o_data_a = 16'b1111110010101000;
            14'h04d7: o_data_a = 16'b1111110000010000;
            14'h04d8: o_data_a = 16'b1110110010100000;
            14'h04d9: o_data_a = 16'b1111000010001000;
            14'h04da: o_data_a = 16'b0000000000000000;
            14'h04db: o_data_a = 16'b1111110010101000;
            14'h04dc: o_data_a = 16'b1111110000010000;
            14'h04dd: o_data_a = 16'b0000000000000011;
            14'h04de: o_data_a = 16'b1111110111100000;
            14'h04df: o_data_a = 16'b1110110111100000;
            14'h04e0: o_data_a = 16'b1110110111100000;
            14'h04e1: o_data_a = 16'b1110110111100000;
            14'h04e2: o_data_a = 16'b1110001100001000;
            14'h04e3: o_data_a = 16'b0000000000000011;
            14'h04e4: o_data_a = 16'b1111110000010000;
            14'h04e5: o_data_a = 16'b0000000000001001;
            14'h04e6: o_data_a = 16'b1110000010100000;
            14'h04e7: o_data_a = 16'b1111110000010000;
            14'h04e8: o_data_a = 16'b0000000000000000;
            14'h04e9: o_data_a = 16'b1111110111101000;
            14'h04ea: o_data_a = 16'b1110110010100000;
            14'h04eb: o_data_a = 16'b1110001100001000;
            14'h04ec: o_data_a = 16'b0000000000000000;
            14'h04ed: o_data_a = 16'b1111110010101000;
            14'h04ee: o_data_a = 16'b1111110000010000;
            14'h04ef: o_data_a = 16'b0000010011110011;
            14'h04f0: o_data_a = 16'b1110001100000101;
            14'h04f1: o_data_a = 16'b0000010100110111;
            14'h04f2: o_data_a = 16'b1110101010000111;
            14'h04f3: o_data_a = 16'b0000000000000011;
            14'h04f4: o_data_a = 16'b1111110000010000;
            14'h04f5: o_data_a = 16'b0000000000000111;
            14'h04f6: o_data_a = 16'b1110000010100000;
            14'h04f7: o_data_a = 16'b1111110000010000;
            14'h04f8: o_data_a = 16'b0000000000000000;
            14'h04f9: o_data_a = 16'b1111110111101000;
            14'h04fa: o_data_a = 16'b1110110010100000;
            14'h04fb: o_data_a = 16'b1110001100001000;
            14'h04fc: o_data_a = 16'b0000000000000000;
            14'h04fd: o_data_a = 16'b1111110010101000;
            14'h04fe: o_data_a = 16'b1111110000010000;
            14'h04ff: o_data_a = 16'b0000010100000011;
            14'h0500: o_data_a = 16'b1110001100000101;
            14'h0501: o_data_a = 16'b0000010100011101;
            14'h0502: o_data_a = 16'b1110101010000111;
            14'h0503: o_data_a = 16'b0000000000000011;
            14'h0504: o_data_a = 16'b1111110000100000;
            14'h0505: o_data_a = 16'b1111110000010000;
            14'h0506: o_data_a = 16'b0000000000000000;
            14'h0507: o_data_a = 16'b1111110111101000;
            14'h0508: o_data_a = 16'b1110110010100000;
            14'h0509: o_data_a = 16'b1110001100001000;
            14'h050a: o_data_a = 16'b0000000000000100;
            14'h050b: o_data_a = 16'b1110110000010000;
            14'h050c: o_data_a = 16'b0000000000000000;
            14'h050d: o_data_a = 16'b1111110111101000;
            14'h050e: o_data_a = 16'b1110110010100000;
            14'h050f: o_data_a = 16'b1110001100001000;
            14'h0510: o_data_a = 16'b0000000000000000;
            14'h0511: o_data_a = 16'b1111110010101000;
            14'h0512: o_data_a = 16'b1111110000010000;
            14'h0513: o_data_a = 16'b1110110010100000;
            14'h0514: o_data_a = 16'b1111000010001000;
            14'h0515: o_data_a = 16'b0000000000000000;
            14'h0516: o_data_a = 16'b1111110010101000;
            14'h0517: o_data_a = 16'b1111110000010000;
            14'h0518: o_data_a = 16'b0000000000000011;
            14'h0519: o_data_a = 16'b1111110000100000;
            14'h051a: o_data_a = 16'b1110001100001000;
            14'h051b: o_data_a = 16'b0000010100110101;
            14'h051c: o_data_a = 16'b1110101010000111;
            14'h051d: o_data_a = 16'b0000000000000011;
            14'h051e: o_data_a = 16'b1111110111100000;
            14'h051f: o_data_a = 16'b1111110000010000;
            14'h0520: o_data_a = 16'b0000000000000000;
            14'h0521: o_data_a = 16'b1111110111101000;
            14'h0522: o_data_a = 16'b1110110010100000;
            14'h0523: o_data_a = 16'b1110001100001000;
            14'h0524: o_data_a = 16'b0000000000000100;
            14'h0525: o_data_a = 16'b1110110000010000;
            14'h0526: o_data_a = 16'b0000000000000000;
            14'h0527: o_data_a = 16'b1111110111101000;
            14'h0528: o_data_a = 16'b1110110010100000;
            14'h0529: o_data_a = 16'b1110001100001000;
            14'h052a: o_data_a = 16'b0000000000000000;
            14'h052b: o_data_a = 16'b1111110010101000;
            14'h052c: o_data_a = 16'b1111110000010000;
            14'h052d: o_data_a = 16'b1110110010100000;
            14'h052e: o_data_a = 16'b1111000010001000;
            14'h052f: o_data_a = 16'b0000000000000000;
            14'h0530: o_data_a = 16'b1111110010101000;
            14'h0531: o_data_a = 16'b1111110000010000;
            14'h0532: o_data_a = 16'b0000000000000011;
            14'h0533: o_data_a = 16'b1111110111100000;
            14'h0534: o_data_a = 16'b1110001100001000;
            14'h0535: o_data_a = 16'b0000010101111001;
            14'h0536: o_data_a = 16'b1110101010000111;
            14'h0537: o_data_a = 16'b0000000000000011;
            14'h0538: o_data_a = 16'b1111110000010000;
            14'h0539: o_data_a = 16'b0000000000000111;
            14'h053a: o_data_a = 16'b1110000010100000;
            14'h053b: o_data_a = 16'b1111110000010000;
            14'h053c: o_data_a = 16'b0000000000000000;
            14'h053d: o_data_a = 16'b1111110111101000;
            14'h053e: o_data_a = 16'b1110110010100000;
            14'h053f: o_data_a = 16'b1110001100001000;
            14'h0540: o_data_a = 16'b0000000000000000;
            14'h0541: o_data_a = 16'b1111110010101000;
            14'h0542: o_data_a = 16'b1111110000010000;
            14'h0543: o_data_a = 16'b0000010101000111;
            14'h0544: o_data_a = 16'b1110001100000101;
            14'h0545: o_data_a = 16'b0000010101100001;
            14'h0546: o_data_a = 16'b1110101010000111;
            14'h0547: o_data_a = 16'b0000000000000011;
            14'h0548: o_data_a = 16'b1111110000100000;
            14'h0549: o_data_a = 16'b1111110000010000;
            14'h054a: o_data_a = 16'b0000000000000000;
            14'h054b: o_data_a = 16'b1111110111101000;
            14'h054c: o_data_a = 16'b1110110010100000;
            14'h054d: o_data_a = 16'b1110001100001000;
            14'h054e: o_data_a = 16'b0000000000000100;
            14'h054f: o_data_a = 16'b1110110000010000;
            14'h0550: o_data_a = 16'b0000000000000000;
            14'h0551: o_data_a = 16'b1111110111101000;
            14'h0552: o_data_a = 16'b1110110010100000;
            14'h0553: o_data_a = 16'b1110001100001000;
            14'h0554: o_data_a = 16'b0000000000000000;
            14'h0555: o_data_a = 16'b1111110010101000;
            14'h0556: o_data_a = 16'b1111110000010000;
            14'h0557: o_data_a = 16'b1110110010100000;
            14'h0558: o_data_a = 16'b1111000111001000;
            14'h0559: o_data_a = 16'b0000000000000000;
            14'h055a: o_data_a = 16'b1111110010101000;
            14'h055b: o_data_a = 16'b1111110000010000;
            14'h055c: o_data_a = 16'b0000000000000011;
            14'h055d: o_data_a = 16'b1111110000100000;
            14'h055e: o_data_a = 16'b1110001100001000;
            14'h055f: o_data_a = 16'b0000010101111001;
            14'h0560: o_data_a = 16'b1110101010000111;
            14'h0561: o_data_a = 16'b0000000000000011;
            14'h0562: o_data_a = 16'b1111110111100000;
            14'h0563: o_data_a = 16'b1111110000010000;
            14'h0564: o_data_a = 16'b0000000000000000;
            14'h0565: o_data_a = 16'b1111110111101000;
            14'h0566: o_data_a = 16'b1110110010100000;
            14'h0567: o_data_a = 16'b1110001100001000;
            14'h0568: o_data_a = 16'b0000000000000100;
            14'h0569: o_data_a = 16'b1110110000010000;
            14'h056a: o_data_a = 16'b0000000000000000;
            14'h056b: o_data_a = 16'b1111110111101000;
            14'h056c: o_data_a = 16'b1110110010100000;
            14'h056d: o_data_a = 16'b1110001100001000;
            14'h056e: o_data_a = 16'b0000000000000000;
            14'h056f: o_data_a = 16'b1111110010101000;
            14'h0570: o_data_a = 16'b1111110000010000;
            14'h0571: o_data_a = 16'b1110110010100000;
            14'h0572: o_data_a = 16'b1111000111001000;
            14'h0573: o_data_a = 16'b0000000000000000;
            14'h0574: o_data_a = 16'b1111110010101000;
            14'h0575: o_data_a = 16'b1111110000010000;
            14'h0576: o_data_a = 16'b0000000000000011;
            14'h0577: o_data_a = 16'b1111110111100000;
            14'h0578: o_data_a = 16'b1110001100001000;
            14'h0579: o_data_a = 16'b0000000000000011;
            14'h057a: o_data_a = 16'b1111110000010000;
            14'h057b: o_data_a = 16'b0000000000001000;
            14'h057c: o_data_a = 16'b1110000010100000;
            14'h057d: o_data_a = 16'b1111110000010000;
            14'h057e: o_data_a = 16'b0000000000000000;
            14'h057f: o_data_a = 16'b1111110111101000;
            14'h0580: o_data_a = 16'b1110110010100000;
            14'h0581: o_data_a = 16'b1110001100001000;
            14'h0582: o_data_a = 16'b0000000000000000;
            14'h0583: o_data_a = 16'b1111110010101000;
            14'h0584: o_data_a = 16'b1111110000010000;
            14'h0585: o_data_a = 16'b0000010110001001;
            14'h0586: o_data_a = 16'b1110001100000101;
            14'h0587: o_data_a = 16'b0000010111001101;
            14'h0588: o_data_a = 16'b1110101010000111;
            14'h0589: o_data_a = 16'b0000000000000011;
            14'h058a: o_data_a = 16'b1111110000010000;
            14'h058b: o_data_a = 16'b0000000000000111;
            14'h058c: o_data_a = 16'b1110000010100000;
            14'h058d: o_data_a = 16'b1111110000010000;
            14'h058e: o_data_a = 16'b0000000000000000;
            14'h058f: o_data_a = 16'b1111110111101000;
            14'h0590: o_data_a = 16'b1110110010100000;
            14'h0591: o_data_a = 16'b1110001100001000;
            14'h0592: o_data_a = 16'b0000000000000000;
            14'h0593: o_data_a = 16'b1111110010101000;
            14'h0594: o_data_a = 16'b1111110000010000;
            14'h0595: o_data_a = 16'b0000010110011001;
            14'h0596: o_data_a = 16'b1110001100000101;
            14'h0597: o_data_a = 16'b0000010110110011;
            14'h0598: o_data_a = 16'b1110101010000111;
            14'h0599: o_data_a = 16'b0000000000000011;
            14'h059a: o_data_a = 16'b1111110111100000;
            14'h059b: o_data_a = 16'b1111110000010000;
            14'h059c: o_data_a = 16'b0000000000000000;
            14'h059d: o_data_a = 16'b1111110111101000;
            14'h059e: o_data_a = 16'b1110110010100000;
            14'h059f: o_data_a = 16'b1110001100001000;
            14'h05a0: o_data_a = 16'b0000000000000100;
            14'h05a1: o_data_a = 16'b1110110000010000;
            14'h05a2: o_data_a = 16'b0000000000000000;
            14'h05a3: o_data_a = 16'b1111110111101000;
            14'h05a4: o_data_a = 16'b1110110010100000;
            14'h05a5: o_data_a = 16'b1110001100001000;
            14'h05a6: o_data_a = 16'b0000000000000000;
            14'h05a7: o_data_a = 16'b1111110010101000;
            14'h05a8: o_data_a = 16'b1111110000010000;
            14'h05a9: o_data_a = 16'b1110110010100000;
            14'h05aa: o_data_a = 16'b1111000010001000;
            14'h05ab: o_data_a = 16'b0000000000000000;
            14'h05ac: o_data_a = 16'b1111110010101000;
            14'h05ad: o_data_a = 16'b1111110000010000;
            14'h05ae: o_data_a = 16'b0000000000000011;
            14'h05af: o_data_a = 16'b1111110111100000;
            14'h05b0: o_data_a = 16'b1110001100001000;
            14'h05b1: o_data_a = 16'b0000010111001011;
            14'h05b2: o_data_a = 16'b1110101010000111;
            14'h05b3: o_data_a = 16'b0000000000000011;
            14'h05b4: o_data_a = 16'b1111110000100000;
            14'h05b5: o_data_a = 16'b1111110000010000;
            14'h05b6: o_data_a = 16'b0000000000000000;
            14'h05b7: o_data_a = 16'b1111110111101000;
            14'h05b8: o_data_a = 16'b1110110010100000;
            14'h05b9: o_data_a = 16'b1110001100001000;
            14'h05ba: o_data_a = 16'b0000000000000100;
            14'h05bb: o_data_a = 16'b1110110000010000;
            14'h05bc: o_data_a = 16'b0000000000000000;
            14'h05bd: o_data_a = 16'b1111110111101000;
            14'h05be: o_data_a = 16'b1110110010100000;
            14'h05bf: o_data_a = 16'b1110001100001000;
            14'h05c0: o_data_a = 16'b0000000000000000;
            14'h05c1: o_data_a = 16'b1111110010101000;
            14'h05c2: o_data_a = 16'b1111110000010000;
            14'h05c3: o_data_a = 16'b1110110010100000;
            14'h05c4: o_data_a = 16'b1111000010001000;
            14'h05c5: o_data_a = 16'b0000000000000000;
            14'h05c6: o_data_a = 16'b1111110010101000;
            14'h05c7: o_data_a = 16'b1111110000010000;
            14'h05c8: o_data_a = 16'b0000000000000011;
            14'h05c9: o_data_a = 16'b1111110000100000;
            14'h05ca: o_data_a = 16'b1110001100001000;
            14'h05cb: o_data_a = 16'b0000011000001111;
            14'h05cc: o_data_a = 16'b1110101010000111;
            14'h05cd: o_data_a = 16'b0000000000000011;
            14'h05ce: o_data_a = 16'b1111110000010000;
            14'h05cf: o_data_a = 16'b0000000000000111;
            14'h05d0: o_data_a = 16'b1110000010100000;
            14'h05d1: o_data_a = 16'b1111110000010000;
            14'h05d2: o_data_a = 16'b0000000000000000;
            14'h05d3: o_data_a = 16'b1111110111101000;
            14'h05d4: o_data_a = 16'b1110110010100000;
            14'h05d5: o_data_a = 16'b1110001100001000;
            14'h05d6: o_data_a = 16'b0000000000000000;
            14'h05d7: o_data_a = 16'b1111110010101000;
            14'h05d8: o_data_a = 16'b1111110000010000;
            14'h05d9: o_data_a = 16'b0000010111011101;
            14'h05da: o_data_a = 16'b1110001100000101;
            14'h05db: o_data_a = 16'b0000010111110111;
            14'h05dc: o_data_a = 16'b1110101010000111;
            14'h05dd: o_data_a = 16'b0000000000000011;
            14'h05de: o_data_a = 16'b1111110111100000;
            14'h05df: o_data_a = 16'b1111110000010000;
            14'h05e0: o_data_a = 16'b0000000000000000;
            14'h05e1: o_data_a = 16'b1111110111101000;
            14'h05e2: o_data_a = 16'b1110110010100000;
            14'h05e3: o_data_a = 16'b1110001100001000;
            14'h05e4: o_data_a = 16'b0000000000000100;
            14'h05e5: o_data_a = 16'b1110110000010000;
            14'h05e6: o_data_a = 16'b0000000000000000;
            14'h05e7: o_data_a = 16'b1111110111101000;
            14'h05e8: o_data_a = 16'b1110110010100000;
            14'h05e9: o_data_a = 16'b1110001100001000;
            14'h05ea: o_data_a = 16'b0000000000000000;
            14'h05eb: o_data_a = 16'b1111110010101000;
            14'h05ec: o_data_a = 16'b1111110000010000;
            14'h05ed: o_data_a = 16'b1110110010100000;
            14'h05ee: o_data_a = 16'b1111000111001000;
            14'h05ef: o_data_a = 16'b0000000000000000;
            14'h05f0: o_data_a = 16'b1111110010101000;
            14'h05f1: o_data_a = 16'b1111110000010000;
            14'h05f2: o_data_a = 16'b0000000000000011;
            14'h05f3: o_data_a = 16'b1111110111100000;
            14'h05f4: o_data_a = 16'b1110001100001000;
            14'h05f5: o_data_a = 16'b0000011000001111;
            14'h05f6: o_data_a = 16'b1110101010000111;
            14'h05f7: o_data_a = 16'b0000000000000011;
            14'h05f8: o_data_a = 16'b1111110000100000;
            14'h05f9: o_data_a = 16'b1111110000010000;
            14'h05fa: o_data_a = 16'b0000000000000000;
            14'h05fb: o_data_a = 16'b1111110111101000;
            14'h05fc: o_data_a = 16'b1110110010100000;
            14'h05fd: o_data_a = 16'b1110001100001000;
            14'h05fe: o_data_a = 16'b0000000000000100;
            14'h05ff: o_data_a = 16'b1110110000010000;
            14'h0600: o_data_a = 16'b0000000000000000;
            14'h0601: o_data_a = 16'b1111110111101000;
            14'h0602: o_data_a = 16'b1110110010100000;
            14'h0603: o_data_a = 16'b1110001100001000;
            14'h0604: o_data_a = 16'b0000000000000000;
            14'h0605: o_data_a = 16'b1111110010101000;
            14'h0606: o_data_a = 16'b1111110000010000;
            14'h0607: o_data_a = 16'b1110110010100000;
            14'h0608: o_data_a = 16'b1111000111001000;
            14'h0609: o_data_a = 16'b0000000000000000;
            14'h060a: o_data_a = 16'b1111110010101000;
            14'h060b: o_data_a = 16'b1111110000010000;
            14'h060c: o_data_a = 16'b0000000000000011;
            14'h060d: o_data_a = 16'b1111110000100000;
            14'h060e: o_data_a = 16'b1110001100001000;
            14'h060f: o_data_a = 16'b0000000000000011;
            14'h0610: o_data_a = 16'b1111110000100000;
            14'h0611: o_data_a = 16'b1111110000010000;
            14'h0612: o_data_a = 16'b0000000000000000;
            14'h0613: o_data_a = 16'b1111110111101000;
            14'h0614: o_data_a = 16'b1110110010100000;
            14'h0615: o_data_a = 16'b1110001100001000;
            14'h0616: o_data_a = 16'b0000000000000011;
            14'h0617: o_data_a = 16'b1111110000010000;
            14'h0618: o_data_a = 16'b0000000000001010;
            14'h0619: o_data_a = 16'b1110000010100000;
            14'h061a: o_data_a = 16'b1111110000010000;
            14'h061b: o_data_a = 16'b0000000000000000;
            14'h061c: o_data_a = 16'b1111110111101000;
            14'h061d: o_data_a = 16'b1110110010100000;
            14'h061e: o_data_a = 16'b1110001100001000;
            14'h061f: o_data_a = 16'b0000011000100011;
            14'h0620: o_data_a = 16'b1110110000010000;
            14'h0621: o_data_a = 16'b0000000000010110;
            14'h0622: o_data_a = 16'b1110101010000111;
            14'h0623: o_data_a = 16'b0000000000000000;
            14'h0624: o_data_a = 16'b1111110010100000;
            14'h0625: o_data_a = 16'b1111110001001000;
            14'h0626: o_data_a = 16'b0000000000000000;
            14'h0627: o_data_a = 16'b1111110010101000;
            14'h0628: o_data_a = 16'b1111110000010000;
            14'h0629: o_data_a = 16'b0000011000101101;
            14'h062a: o_data_a = 16'b1110001100000101;
            14'h062b: o_data_a = 16'b0000011001001100;
            14'h062c: o_data_a = 16'b1110101010000111;
            14'h062d: o_data_a = 16'b0000000000000000;
            14'h062e: o_data_a = 16'b1111110111001000;
            14'h062f: o_data_a = 16'b1111110010100000;
            14'h0630: o_data_a = 16'b1110111111001000;
            14'h0631: o_data_a = 16'b0000000000000011;
            14'h0632: o_data_a = 16'b1111110000010000;
            14'h0633: o_data_a = 16'b0000000000001110;
            14'h0634: o_data_a = 16'b1110000010010000;
            14'h0635: o_data_a = 16'b0000000000001101;
            14'h0636: o_data_a = 16'b1110001100001000;
            14'h0637: o_data_a = 16'b0000000000000000;
            14'h0638: o_data_a = 16'b1111110010101000;
            14'h0639: o_data_a = 16'b1111110000010000;
            14'h063a: o_data_a = 16'b0000000000001101;
            14'h063b: o_data_a = 16'b1111110000100000;
            14'h063c: o_data_a = 16'b1110001100001000;
            14'h063d: o_data_a = 16'b0000000000000011;
            14'h063e: o_data_a = 16'b1111110000010000;
            14'h063f: o_data_a = 16'b0000000000001010;
            14'h0640: o_data_a = 16'b1110000010100000;
            14'h0641: o_data_a = 16'b1111110000010000;
            14'h0642: o_data_a = 16'b0000000000000000;
            14'h0643: o_data_a = 16'b1111110111101000;
            14'h0644: o_data_a = 16'b1110110010100000;
            14'h0645: o_data_a = 16'b1110001100001000;
            14'h0646: o_data_a = 16'b0000000000000000;
            14'h0647: o_data_a = 16'b1111110010101000;
            14'h0648: o_data_a = 16'b1111110000010000;
            14'h0649: o_data_a = 16'b0000000000000011;
            14'h064a: o_data_a = 16'b1111110000100000;
            14'h064b: o_data_a = 16'b1110001100001000;
            14'h064c: o_data_a = 16'b0000000000000011;
            14'h064d: o_data_a = 16'b1111110000100000;
            14'h064e: o_data_a = 16'b1111110000010000;
            14'h064f: o_data_a = 16'b0000000000000000;
            14'h0650: o_data_a = 16'b1111110111101000;
            14'h0651: o_data_a = 16'b1110110010100000;
            14'h0652: o_data_a = 16'b1110001100001000;
            14'h0653: o_data_a = 16'b0000000000000011;
            14'h0654: o_data_a = 16'b1111110000010000;
            14'h0655: o_data_a = 16'b0000000000001011;
            14'h0656: o_data_a = 16'b1110000010100000;
            14'h0657: o_data_a = 16'b1111110000010000;
            14'h0658: o_data_a = 16'b0000000000000000;
            14'h0659: o_data_a = 16'b1111110111101000;
            14'h065a: o_data_a = 16'b1110110010100000;
            14'h065b: o_data_a = 16'b1110001100001000;
            14'h065c: o_data_a = 16'b0000011001100000;
            14'h065d: o_data_a = 16'b1110110000010000;
            14'h065e: o_data_a = 16'b0000000000100110;
            14'h065f: o_data_a = 16'b1110101010000111;
            14'h0660: o_data_a = 16'b0000000000000000;
            14'h0661: o_data_a = 16'b1111110010100000;
            14'h0662: o_data_a = 16'b1111110001001000;
            14'h0663: o_data_a = 16'b0000000000000000;
            14'h0664: o_data_a = 16'b1111110010101000;
            14'h0665: o_data_a = 16'b1111110000010000;
            14'h0666: o_data_a = 16'b0000011001101010;
            14'h0667: o_data_a = 16'b1110001100000101;
            14'h0668: o_data_a = 16'b0000011010001011;
            14'h0669: o_data_a = 16'b1110101010000111;
            14'h066a: o_data_a = 16'b0000000000000010;
            14'h066b: o_data_a = 16'b1110110000010000;
            14'h066c: o_data_a = 16'b0000000000000000;
            14'h066d: o_data_a = 16'b1111110111101000;
            14'h066e: o_data_a = 16'b1110110010100000;
            14'h066f: o_data_a = 16'b1110001100001000;
            14'h0670: o_data_a = 16'b0000000000000011;
            14'h0671: o_data_a = 16'b1111110000010000;
            14'h0672: o_data_a = 16'b0000000000001110;
            14'h0673: o_data_a = 16'b1110000010010000;
            14'h0674: o_data_a = 16'b0000000000001101;
            14'h0675: o_data_a = 16'b1110001100001000;
            14'h0676: o_data_a = 16'b0000000000000000;
            14'h0677: o_data_a = 16'b1111110010101000;
            14'h0678: o_data_a = 16'b1111110000010000;
            14'h0679: o_data_a = 16'b0000000000001101;
            14'h067a: o_data_a = 16'b1111110000100000;
            14'h067b: o_data_a = 16'b1110001100001000;
            14'h067c: o_data_a = 16'b0000000000000011;
            14'h067d: o_data_a = 16'b1111110000010000;
            14'h067e: o_data_a = 16'b0000000000001011;
            14'h067f: o_data_a = 16'b1110000010100000;
            14'h0680: o_data_a = 16'b1111110000010000;
            14'h0681: o_data_a = 16'b0000000000000000;
            14'h0682: o_data_a = 16'b1111110111101000;
            14'h0683: o_data_a = 16'b1110110010100000;
            14'h0684: o_data_a = 16'b1110001100001000;
            14'h0685: o_data_a = 16'b0000000000000000;
            14'h0686: o_data_a = 16'b1111110010101000;
            14'h0687: o_data_a = 16'b1111110000010000;
            14'h0688: o_data_a = 16'b0000000000000011;
            14'h0689: o_data_a = 16'b1111110000100000;
            14'h068a: o_data_a = 16'b1110001100001000;
            14'h068b: o_data_a = 16'b0000000000000011;
            14'h068c: o_data_a = 16'b1111110111100000;
            14'h068d: o_data_a = 16'b1111110000010000;
            14'h068e: o_data_a = 16'b0000000000000000;
            14'h068f: o_data_a = 16'b1111110111101000;
            14'h0690: o_data_a = 16'b1110110010100000;
            14'h0691: o_data_a = 16'b1110001100001000;
            14'h0692: o_data_a = 16'b0000000000000011;
            14'h0693: o_data_a = 16'b1111110000010000;
            14'h0694: o_data_a = 16'b0000000000001100;
            14'h0695: o_data_a = 16'b1110000010100000;
            14'h0696: o_data_a = 16'b1111110000010000;
            14'h0697: o_data_a = 16'b0000000000000000;
            14'h0698: o_data_a = 16'b1111110111101000;
            14'h0699: o_data_a = 16'b1110110010100000;
            14'h069a: o_data_a = 16'b1110001100001000;
            14'h069b: o_data_a = 16'b0000011010011111;
            14'h069c: o_data_a = 16'b1110110000010000;
            14'h069d: o_data_a = 16'b0000000000010110;
            14'h069e: o_data_a = 16'b1110101010000111;
            14'h069f: o_data_a = 16'b0000000000000000;
            14'h06a0: o_data_a = 16'b1111110010100000;
            14'h06a1: o_data_a = 16'b1111110001001000;
            14'h06a2: o_data_a = 16'b0000000000000000;
            14'h06a3: o_data_a = 16'b1111110010101000;
            14'h06a4: o_data_a = 16'b1111110000010000;
            14'h06a5: o_data_a = 16'b0000011010101001;
            14'h06a6: o_data_a = 16'b1110001100000101;
            14'h06a7: o_data_a = 16'b0000011011001010;
            14'h06a8: o_data_a = 16'b1110101010000111;
            14'h06a9: o_data_a = 16'b0000000000000011;
            14'h06aa: o_data_a = 16'b1110110000010000;
            14'h06ab: o_data_a = 16'b0000000000000000;
            14'h06ac: o_data_a = 16'b1111110111101000;
            14'h06ad: o_data_a = 16'b1110110010100000;
            14'h06ae: o_data_a = 16'b1110001100001000;
            14'h06af: o_data_a = 16'b0000000000000011;
            14'h06b0: o_data_a = 16'b1111110000010000;
            14'h06b1: o_data_a = 16'b0000000000001110;
            14'h06b2: o_data_a = 16'b1110000010010000;
            14'h06b3: o_data_a = 16'b0000000000001101;
            14'h06b4: o_data_a = 16'b1110001100001000;
            14'h06b5: o_data_a = 16'b0000000000000000;
            14'h06b6: o_data_a = 16'b1111110010101000;
            14'h06b7: o_data_a = 16'b1111110000010000;
            14'h06b8: o_data_a = 16'b0000000000001101;
            14'h06b9: o_data_a = 16'b1111110000100000;
            14'h06ba: o_data_a = 16'b1110001100001000;
            14'h06bb: o_data_a = 16'b0000000000000011;
            14'h06bc: o_data_a = 16'b1111110000010000;
            14'h06bd: o_data_a = 16'b0000000000001100;
            14'h06be: o_data_a = 16'b1110000010100000;
            14'h06bf: o_data_a = 16'b1111110000010000;
            14'h06c0: o_data_a = 16'b0000000000000000;
            14'h06c1: o_data_a = 16'b1111110111101000;
            14'h06c2: o_data_a = 16'b1110110010100000;
            14'h06c3: o_data_a = 16'b1110001100001000;
            14'h06c4: o_data_a = 16'b0000000000000000;
            14'h06c5: o_data_a = 16'b1111110010101000;
            14'h06c6: o_data_a = 16'b1111110000010000;
            14'h06c7: o_data_a = 16'b0000000000000011;
            14'h06c8: o_data_a = 16'b1111110111100000;
            14'h06c9: o_data_a = 16'b1110001100001000;
            14'h06ca: o_data_a = 16'b0000000000000011;
            14'h06cb: o_data_a = 16'b1111110111100000;
            14'h06cc: o_data_a = 16'b1111110000010000;
            14'h06cd: o_data_a = 16'b0000000000000000;
            14'h06ce: o_data_a = 16'b1111110111101000;
            14'h06cf: o_data_a = 16'b1110110010100000;
            14'h06d0: o_data_a = 16'b1110001100001000;
            14'h06d1: o_data_a = 16'b0000000000000011;
            14'h06d2: o_data_a = 16'b1111110000010000;
            14'h06d3: o_data_a = 16'b0000000000001101;
            14'h06d4: o_data_a = 16'b1110000010100000;
            14'h06d5: o_data_a = 16'b1111110000010000;
            14'h06d6: o_data_a = 16'b0000000000000000;
            14'h06d7: o_data_a = 16'b1111110111101000;
            14'h06d8: o_data_a = 16'b1110110010100000;
            14'h06d9: o_data_a = 16'b1110001100001000;
            14'h06da: o_data_a = 16'b0000011011011110;
            14'h06db: o_data_a = 16'b1110110000010000;
            14'h06dc: o_data_a = 16'b0000000000100110;
            14'h06dd: o_data_a = 16'b1110101010000111;
            14'h06de: o_data_a = 16'b0000000000000000;
            14'h06df: o_data_a = 16'b1111110010100000;
            14'h06e0: o_data_a = 16'b1111110001001000;
            14'h06e1: o_data_a = 16'b0000000000000000;
            14'h06e2: o_data_a = 16'b1111110010101000;
            14'h06e3: o_data_a = 16'b1111110000010000;
            14'h06e4: o_data_a = 16'b0000011011101000;
            14'h06e5: o_data_a = 16'b1110001100000101;
            14'h06e6: o_data_a = 16'b0000011100001001;
            14'h06e7: o_data_a = 16'b1110101010000111;
            14'h06e8: o_data_a = 16'b0000000000000100;
            14'h06e9: o_data_a = 16'b1110110000010000;
            14'h06ea: o_data_a = 16'b0000000000000000;
            14'h06eb: o_data_a = 16'b1111110111101000;
            14'h06ec: o_data_a = 16'b1110110010100000;
            14'h06ed: o_data_a = 16'b1110001100001000;
            14'h06ee: o_data_a = 16'b0000000000000011;
            14'h06ef: o_data_a = 16'b1111110000010000;
            14'h06f0: o_data_a = 16'b0000000000001110;
            14'h06f1: o_data_a = 16'b1110000010010000;
            14'h06f2: o_data_a = 16'b0000000000001101;
            14'h06f3: o_data_a = 16'b1110001100001000;
            14'h06f4: o_data_a = 16'b0000000000000000;
            14'h06f5: o_data_a = 16'b1111110010101000;
            14'h06f6: o_data_a = 16'b1111110000010000;
            14'h06f7: o_data_a = 16'b0000000000001101;
            14'h06f8: o_data_a = 16'b1111110000100000;
            14'h06f9: o_data_a = 16'b1110001100001000;
            14'h06fa: o_data_a = 16'b0000000000000011;
            14'h06fb: o_data_a = 16'b1111110000010000;
            14'h06fc: o_data_a = 16'b0000000000001101;
            14'h06fd: o_data_a = 16'b1110000010100000;
            14'h06fe: o_data_a = 16'b1111110000010000;
            14'h06ff: o_data_a = 16'b0000000000000000;
            14'h0700: o_data_a = 16'b1111110111101000;
            14'h0701: o_data_a = 16'b1110110010100000;
            14'h0702: o_data_a = 16'b1110001100001000;
            14'h0703: o_data_a = 16'b0000000000000000;
            14'h0704: o_data_a = 16'b1111110010101000;
            14'h0705: o_data_a = 16'b1111110000010000;
            14'h0706: o_data_a = 16'b0000000000000011;
            14'h0707: o_data_a = 16'b1111110111100000;
            14'h0708: o_data_a = 16'b1110001100001000;
            14'h0709: o_data_a = 16'b0000000000000011;
            14'h070a: o_data_a = 16'b1111110000010000;
            14'h070b: o_data_a = 16'b0000000000000000;
            14'h070c: o_data_a = 16'b1111110111101000;
            14'h070d: o_data_a = 16'b1110110010100000;
            14'h070e: o_data_a = 16'b1110001100001000;
            14'h070f: o_data_a = 16'b0000000000000001;
            14'h0710: o_data_a = 16'b1110110000010000;
            14'h0711: o_data_a = 16'b0000000000001101;
            14'h0712: o_data_a = 16'b1110001100001000;
            14'h0713: o_data_a = 16'b0000000110000011;
            14'h0714: o_data_a = 16'b1110110000010000;
            14'h0715: o_data_a = 16'b0000000000001110;
            14'h0716: o_data_a = 16'b1110001100001000;
            14'h0717: o_data_a = 16'b0000011100011011;
            14'h0718: o_data_a = 16'b1110110000010000;
            14'h0719: o_data_a = 16'b0000000001011111;
            14'h071a: o_data_a = 16'b1110101010000111;
            14'h071b: o_data_a = 16'b0000000000000000;
            14'h071c: o_data_a = 16'b1111110010101000;
            14'h071d: o_data_a = 16'b1111110000010000;
            14'h071e: o_data_a = 16'b0000000000000101;
            14'h071f: o_data_a = 16'b1110001100001000;
            14'h0720: o_data_a = 16'b0000000000000011;
            14'h0721: o_data_a = 16'b1111110000010000;
            14'h0722: o_data_a = 16'b0000000000001110;
            14'h0723: o_data_a = 16'b1110000010100000;
            14'h0724: o_data_a = 16'b1111110000010000;
            14'h0725: o_data_a = 16'b0000000000000000;
            14'h0726: o_data_a = 16'b1111110111101000;
            14'h0727: o_data_a = 16'b1110110010100000;
            14'h0728: o_data_a = 16'b1110001100001000;
            14'h0729: o_data_a = 16'b0000000000110110;
            14'h072a: o_data_a = 16'b1110101010000111;
            14'h072b: o_data_a = 16'b0000000000000101;
            14'h072c: o_data_a = 16'b1110110000010000;
            14'h072d: o_data_a = 16'b1110001110010000;
            14'h072e: o_data_a = 16'b0000000000000000;
            14'h072f: o_data_a = 16'b1111110111101000;
            14'h0730: o_data_a = 16'b1110110010100000;
            14'h0731: o_data_a = 16'b1110101010001000;
            14'h0732: o_data_a = 16'b0000011100101101;
            14'h0733: o_data_a = 16'b1110001100000001;
            14'h0734: o_data_a = 16'b0000000000000010;
            14'h0735: o_data_a = 16'b1111110000100000;
            14'h0736: o_data_a = 16'b1111110000010000;
            14'h0737: o_data_a = 16'b0000000000000000;
            14'h0738: o_data_a = 16'b1111110111101000;
            14'h0739: o_data_a = 16'b1110110010100000;
            14'h073a: o_data_a = 16'b1110001100001000;
            14'h073b: o_data_a = 16'b0000000000000000;
            14'h073c: o_data_a = 16'b1111110010101000;
            14'h073d: o_data_a = 16'b1111110000010000;
            14'h073e: o_data_a = 16'b0000000000000011;
            14'h073f: o_data_a = 16'b1110001100001000;
            14'h0740: o_data_a = 16'b0000000000000011;
            14'h0741: o_data_a = 16'b1111110111100000;
            14'h0742: o_data_a = 16'b1110110111100000;
            14'h0743: o_data_a = 16'b1111110000010000;
            14'h0744: o_data_a = 16'b0000000000000000;
            14'h0745: o_data_a = 16'b1111110111101000;
            14'h0746: o_data_a = 16'b1110110010100000;
            14'h0747: o_data_a = 16'b1110001100001000;
            14'h0748: o_data_a = 16'b0000000000001010;
            14'h0749: o_data_a = 16'b1110110000010000;
            14'h074a: o_data_a = 16'b0000000000000000;
            14'h074b: o_data_a = 16'b1111110111101000;
            14'h074c: o_data_a = 16'b1110110010100000;
            14'h074d: o_data_a = 16'b1110001100001000;
            14'h074e: o_data_a = 16'b0000000000000010;
            14'h074f: o_data_a = 16'b1110110000010000;
            14'h0750: o_data_a = 16'b0000000000001101;
            14'h0751: o_data_a = 16'b1110001100001000;
            14'h0752: o_data_a = 16'b0001110001110111;
            14'h0753: o_data_a = 16'b1110110000010000;
            14'h0754: o_data_a = 16'b0000000000001110;
            14'h0755: o_data_a = 16'b1110001100001000;
            14'h0756: o_data_a = 16'b0000011101011010;
            14'h0757: o_data_a = 16'b1110110000010000;
            14'h0758: o_data_a = 16'b0000000001011111;
            14'h0759: o_data_a = 16'b1110101010000111;
            14'h075a: o_data_a = 16'b0000000000000000;
            14'h075b: o_data_a = 16'b1111110010101000;
            14'h075c: o_data_a = 16'b1111110000010000;
            14'h075d: o_data_a = 16'b0000000000000001;
            14'h075e: o_data_a = 16'b1111110111100000;
            14'h075f: o_data_a = 16'b1110110111100000;
            14'h0760: o_data_a = 16'b1110001100001000;
            14'h0761: o_data_a = 16'b0000000000000011;
            14'h0762: o_data_a = 16'b1111110000010000;
            14'h0763: o_data_a = 16'b0000000000000011;
            14'h0764: o_data_a = 16'b1110000010100000;
            14'h0765: o_data_a = 16'b1111110000010000;
            14'h0766: o_data_a = 16'b0000000000000000;
            14'h0767: o_data_a = 16'b1111110111101000;
            14'h0768: o_data_a = 16'b1110110010100000;
            14'h0769: o_data_a = 16'b1110001100001000;
            14'h076a: o_data_a = 16'b0000000000001010;
            14'h076b: o_data_a = 16'b1110110000010000;
            14'h076c: o_data_a = 16'b0000000000000000;
            14'h076d: o_data_a = 16'b1111110111101000;
            14'h076e: o_data_a = 16'b1110110010100000;
            14'h076f: o_data_a = 16'b1110001100001000;
            14'h0770: o_data_a = 16'b0000000000000010;
            14'h0771: o_data_a = 16'b1110110000010000;
            14'h0772: o_data_a = 16'b0000000000001101;
            14'h0773: o_data_a = 16'b1110001100001000;
            14'h0774: o_data_a = 16'b0001110001110111;
            14'h0775: o_data_a = 16'b1110110000010000;
            14'h0776: o_data_a = 16'b0000000000001110;
            14'h0777: o_data_a = 16'b1110001100001000;
            14'h0778: o_data_a = 16'b0000011101111100;
            14'h0779: o_data_a = 16'b1110110000010000;
            14'h077a: o_data_a = 16'b0000000001011111;
            14'h077b: o_data_a = 16'b1110101010000111;
            14'h077c: o_data_a = 16'b0000000000000000;
            14'h077d: o_data_a = 16'b1111110010101000;
            14'h077e: o_data_a = 16'b1111110000010000;
            14'h077f: o_data_a = 16'b0000000000000001;
            14'h0780: o_data_a = 16'b1111110111100000;
            14'h0781: o_data_a = 16'b1110110111100000;
            14'h0782: o_data_a = 16'b1110110111100000;
            14'h0783: o_data_a = 16'b1110001100001000;
            14'h0784: o_data_a = 16'b0000000000000010;
            14'h0785: o_data_a = 16'b1111110111100000;
            14'h0786: o_data_a = 16'b1111110000010000;
            14'h0787: o_data_a = 16'b0000000000000000;
            14'h0788: o_data_a = 16'b1111110111101000;
            14'h0789: o_data_a = 16'b1110110010100000;
            14'h078a: o_data_a = 16'b1110001100001000;
            14'h078b: o_data_a = 16'b0000000000000000;
            14'h078c: o_data_a = 16'b1111110111001000;
            14'h078d: o_data_a = 16'b1111110010100000;
            14'h078e: o_data_a = 16'b1110101010001000;
            14'h078f: o_data_a = 16'b0000011110010011;
            14'h0790: o_data_a = 16'b1110110000010000;
            14'h0791: o_data_a = 16'b0000000000000110;
            14'h0792: o_data_a = 16'b1110101010000111;
            14'h0793: o_data_a = 16'b0000000000000000;
            14'h0794: o_data_a = 16'b1111110010101000;
            14'h0795: o_data_a = 16'b1111110000010000;
            14'h0796: o_data_a = 16'b0000011110011010;
            14'h0797: o_data_a = 16'b1110001100000101;
            14'h0798: o_data_a = 16'b0000011110101011;
            14'h0799: o_data_a = 16'b1110101010000111;
            14'h079a: o_data_a = 16'b0000000000001010;
            14'h079b: o_data_a = 16'b1110110000010000;
            14'h079c: o_data_a = 16'b0000000000000000;
            14'h079d: o_data_a = 16'b1111110111101000;
            14'h079e: o_data_a = 16'b1110110010100000;
            14'h079f: o_data_a = 16'b1110001100001000;
            14'h07a0: o_data_a = 16'b0000000000000000;
            14'h07a1: o_data_a = 16'b1111110010101000;
            14'h07a2: o_data_a = 16'b1111110000010000;
            14'h07a3: o_data_a = 16'b0000000000000001;
            14'h07a4: o_data_a = 16'b1111110111100000;
            14'h07a5: o_data_a = 16'b1110110111100000;
            14'h07a6: o_data_a = 16'b1110110111100000;
            14'h07a7: o_data_a = 16'b1110110111100000;
            14'h07a8: o_data_a = 16'b1110001100001000;
            14'h07a9: o_data_a = 16'b0000100000100110;
            14'h07aa: o_data_a = 16'b1110101010000111;
            14'h07ab: o_data_a = 16'b0000000000000011;
            14'h07ac: o_data_a = 16'b1111110111100000;
            14'h07ad: o_data_a = 16'b1110110111100000;
            14'h07ae: o_data_a = 16'b1111110000010000;
            14'h07af: o_data_a = 16'b0000000000000000;
            14'h07b0: o_data_a = 16'b1111110111101000;
            14'h07b1: o_data_a = 16'b1110110010100000;
            14'h07b2: o_data_a = 16'b1110001100001000;
            14'h07b3: o_data_a = 16'b0000000000000000;
            14'h07b4: o_data_a = 16'b1111110111001000;
            14'h07b5: o_data_a = 16'b1111110010100000;
            14'h07b6: o_data_a = 16'b1110101010001000;
            14'h07b7: o_data_a = 16'b0000011110111011;
            14'h07b8: o_data_a = 16'b1110110000010000;
            14'h07b9: o_data_a = 16'b0000000000100110;
            14'h07ba: o_data_a = 16'b1110101010000111;
            14'h07bb: o_data_a = 16'b0000000000000000;
            14'h07bc: o_data_a = 16'b1111110010100000;
            14'h07bd: o_data_a = 16'b1111110001001000;
            14'h07be: o_data_a = 16'b0000000000000010;
            14'h07bf: o_data_a = 16'b1111110111100000;
            14'h07c0: o_data_a = 16'b1111110000010000;
            14'h07c1: o_data_a = 16'b0000000000000000;
            14'h07c2: o_data_a = 16'b1111110111101000;
            14'h07c3: o_data_a = 16'b1110110010100000;
            14'h07c4: o_data_a = 16'b1110001100001000;
            14'h07c5: o_data_a = 16'b0000000000000000;
            14'h07c6: o_data_a = 16'b1111110111001000;
            14'h07c7: o_data_a = 16'b1111110010100000;
            14'h07c8: o_data_a = 16'b1110111111001000;
            14'h07c9: o_data_a = 16'b0000011111001101;
            14'h07ca: o_data_a = 16'b1110110000010000;
            14'h07cb: o_data_a = 16'b0000000000000110;
            14'h07cc: o_data_a = 16'b1110101010000111;
            14'h07cd: o_data_a = 16'b0000000000000000;
            14'h07ce: o_data_a = 16'b1111110010101000;
            14'h07cf: o_data_a = 16'b1111110000010000;
            14'h07d0: o_data_a = 16'b1110110010100000;
            14'h07d1: o_data_a = 16'b1111000000001000;
            14'h07d2: o_data_a = 16'b0000000000000011;
            14'h07d3: o_data_a = 16'b1111110111100000;
            14'h07d4: o_data_a = 16'b1110110111100000;
            14'h07d5: o_data_a = 16'b1111110000010000;
            14'h07d6: o_data_a = 16'b0000000000000000;
            14'h07d7: o_data_a = 16'b1111110111101000;
            14'h07d8: o_data_a = 16'b1110110010100000;
            14'h07d9: o_data_a = 16'b1110001100001000;
            14'h07da: o_data_a = 16'b0000000000000000;
            14'h07db: o_data_a = 16'b1111110111001000;
            14'h07dc: o_data_a = 16'b1111110010100000;
            14'h07dd: o_data_a = 16'b1110101010001000;
            14'h07de: o_data_a = 16'b0000011111100010;
            14'h07df: o_data_a = 16'b1110110000010000;
            14'h07e0: o_data_a = 16'b0000000000100110;
            14'h07e1: o_data_a = 16'b1110101010000111;
            14'h07e2: o_data_a = 16'b0000000000000000;
            14'h07e3: o_data_a = 16'b1111110010101000;
            14'h07e4: o_data_a = 16'b1111110000010000;
            14'h07e5: o_data_a = 16'b1110110010100000;
            14'h07e6: o_data_a = 16'b1111010101001000;
            14'h07e7: o_data_a = 16'b0000000000000010;
            14'h07e8: o_data_a = 16'b1111110111100000;
            14'h07e9: o_data_a = 16'b1111110000010000;
            14'h07ea: o_data_a = 16'b0000000000000000;
            14'h07eb: o_data_a = 16'b1111110111101000;
            14'h07ec: o_data_a = 16'b1110110010100000;
            14'h07ed: o_data_a = 16'b1110001100001000;
            14'h07ee: o_data_a = 16'b0000000000000000;
            14'h07ef: o_data_a = 16'b1111110111001000;
            14'h07f0: o_data_a = 16'b1111110010100000;
            14'h07f1: o_data_a = 16'b1110111111001000;
            14'h07f2: o_data_a = 16'b0000000000000000;
            14'h07f3: o_data_a = 16'b1111110010100000;
            14'h07f4: o_data_a = 16'b1111110001010000;
            14'h07f5: o_data_a = 16'b1110011111001000;
            14'h07f6: o_data_a = 16'b0000011111111010;
            14'h07f7: o_data_a = 16'b1110110000010000;
            14'h07f8: o_data_a = 16'b0000000000000110;
            14'h07f9: o_data_a = 16'b1110101010000111;
            14'h07fa: o_data_a = 16'b0000000000000000;
            14'h07fb: o_data_a = 16'b1111110010101000;
            14'h07fc: o_data_a = 16'b1111110000010000;
            14'h07fd: o_data_a = 16'b1110110010100000;
            14'h07fe: o_data_a = 16'b1111000000001000;
            14'h07ff: o_data_a = 16'b0000000000000000;
            14'h0800: o_data_a = 16'b1111110010101000;
            14'h0801: o_data_a = 16'b1111110000010000;
            14'h0802: o_data_a = 16'b0000100000000110;
            14'h0803: o_data_a = 16'b1110001100000101;
            14'h0804: o_data_a = 16'b0000100000010111;
            14'h0805: o_data_a = 16'b1110101010000111;
            14'h0806: o_data_a = 16'b0000000000010100;
            14'h0807: o_data_a = 16'b1110110000010000;
            14'h0808: o_data_a = 16'b0000000000000000;
            14'h0809: o_data_a = 16'b1111110111101000;
            14'h080a: o_data_a = 16'b1110110010100000;
            14'h080b: o_data_a = 16'b1110001100001000;
            14'h080c: o_data_a = 16'b0000000000000000;
            14'h080d: o_data_a = 16'b1111110010101000;
            14'h080e: o_data_a = 16'b1111110000010000;
            14'h080f: o_data_a = 16'b0000000000000001;
            14'h0810: o_data_a = 16'b1111110111100000;
            14'h0811: o_data_a = 16'b1110110111100000;
            14'h0812: o_data_a = 16'b1110110111100000;
            14'h0813: o_data_a = 16'b1110110111100000;
            14'h0814: o_data_a = 16'b1110001100001000;
            14'h0815: o_data_a = 16'b0000100000100110;
            14'h0816: o_data_a = 16'b1110101010000111;
            14'h0817: o_data_a = 16'b0000000000000101;
            14'h0818: o_data_a = 16'b1110110000010000;
            14'h0819: o_data_a = 16'b0000000000000000;
            14'h081a: o_data_a = 16'b1111110111101000;
            14'h081b: o_data_a = 16'b1110110010100000;
            14'h081c: o_data_a = 16'b1110001100001000;
            14'h081d: o_data_a = 16'b0000000000000000;
            14'h081e: o_data_a = 16'b1111110010101000;
            14'h081f: o_data_a = 16'b1111110000010000;
            14'h0820: o_data_a = 16'b0000000000000001;
            14'h0821: o_data_a = 16'b1111110111100000;
            14'h0822: o_data_a = 16'b1110110111100000;
            14'h0823: o_data_a = 16'b1110110111100000;
            14'h0824: o_data_a = 16'b1110110111100000;
            14'h0825: o_data_a = 16'b1110001100001000;
            14'h0826: o_data_a = 16'b0000000000000011;
            14'h0827: o_data_a = 16'b1111110000010000;
            14'h0828: o_data_a = 16'b0000000000001110;
            14'h0829: o_data_a = 16'b1110000010100000;
            14'h082a: o_data_a = 16'b1111110000010000;
            14'h082b: o_data_a = 16'b0000000000000000;
            14'h082c: o_data_a = 16'b1111110111101000;
            14'h082d: o_data_a = 16'b1110110010100000;
            14'h082e: o_data_a = 16'b1110001100001000;
            14'h082f: o_data_a = 16'b0000000000000000;
            14'h0830: o_data_a = 16'b1111110111001000;
            14'h0831: o_data_a = 16'b1111110010100000;
            14'h0832: o_data_a = 16'b1110111111001000;
            14'h0833: o_data_a = 16'b0000100000110111;
            14'h0834: o_data_a = 16'b1110110000010000;
            14'h0835: o_data_a = 16'b0000000000000110;
            14'h0836: o_data_a = 16'b1110101010000111;
            14'h0837: o_data_a = 16'b0000000000000000;
            14'h0838: o_data_a = 16'b1111110010101000;
            14'h0839: o_data_a = 16'b1111110000010000;
            14'h083a: o_data_a = 16'b0000100000111110;
            14'h083b: o_data_a = 16'b1110001100000101;
            14'h083c: o_data_a = 16'b0000100010110011;
            14'h083d: o_data_a = 16'b1110101010000111;
            14'h083e: o_data_a = 16'b0000000111111010;
            14'h083f: o_data_a = 16'b1110110000010000;
            14'h0840: o_data_a = 16'b0000000000000000;
            14'h0841: o_data_a = 16'b1111110111101000;
            14'h0842: o_data_a = 16'b1110110010100000;
            14'h0843: o_data_a = 16'b1110001100001000;
            14'h0844: o_data_a = 16'b0000000000000000;
            14'h0845: o_data_a = 16'b1111110010101000;
            14'h0846: o_data_a = 16'b1111110000010000;
            14'h0847: o_data_a = 16'b0000000000000001;
            14'h0848: o_data_a = 16'b1111110000100000;
            14'h0849: o_data_a = 16'b1110001100001000;
            14'h084a: o_data_a = 16'b0000000000000001;
            14'h084b: o_data_a = 16'b1111110000010000;
            14'h084c: o_data_a = 16'b0000000000000011;
            14'h084d: o_data_a = 16'b1110000010100000;
            14'h084e: o_data_a = 16'b1111110000010000;
            14'h084f: o_data_a = 16'b0000000000000000;
            14'h0850: o_data_a = 16'b1111110111101000;
            14'h0851: o_data_a = 16'b1110110010100000;
            14'h0852: o_data_a = 16'b1110001100001000;
            14'h0853: o_data_a = 16'b0000000000110010;
            14'h0854: o_data_a = 16'b1110110000010000;
            14'h0855: o_data_a = 16'b0000000000000000;
            14'h0856: o_data_a = 16'b1111110111101000;
            14'h0857: o_data_a = 16'b1110110010100000;
            14'h0858: o_data_a = 16'b1110001100001000;
            14'h0859: o_data_a = 16'b0000000000000000;
            14'h085a: o_data_a = 16'b1111110010100000;
            14'h085b: o_data_a = 16'b1111110001010000;
            14'h085c: o_data_a = 16'b1110011111001000;
            14'h085d: o_data_a = 16'b0000000000000010;
            14'h085e: o_data_a = 16'b1110110000010000;
            14'h085f: o_data_a = 16'b0000000000001101;
            14'h0860: o_data_a = 16'b1110001100001000;
            14'h0861: o_data_a = 16'b0001101010100110;
            14'h0862: o_data_a = 16'b1110110000010000;
            14'h0863: o_data_a = 16'b0000000000001110;
            14'h0864: o_data_a = 16'b1110001100001000;
            14'h0865: o_data_a = 16'b0000100001101001;
            14'h0866: o_data_a = 16'b1110110000010000;
            14'h0867: o_data_a = 16'b0000000001011111;
            14'h0868: o_data_a = 16'b1110101010000111;
            14'h0869: o_data_a = 16'b0000000000000001;
            14'h086a: o_data_a = 16'b1111110111100000;
            14'h086b: o_data_a = 16'b1110110111100000;
            14'h086c: o_data_a = 16'b1111110000010000;
            14'h086d: o_data_a = 16'b0000000000000000;
            14'h086e: o_data_a = 16'b1111110111101000;
            14'h086f: o_data_a = 16'b1110110010100000;
            14'h0870: o_data_a = 16'b1110001100001000;
            14'h0871: o_data_a = 16'b0000000000000010;
            14'h0872: o_data_a = 16'b1110110000010000;
            14'h0873: o_data_a = 16'b0000000000001101;
            14'h0874: o_data_a = 16'b1110001100001000;
            14'h0875: o_data_a = 16'b0001110001110111;
            14'h0876: o_data_a = 16'b1110110000010000;
            14'h0877: o_data_a = 16'b0000000000001110;
            14'h0878: o_data_a = 16'b1110001100001000;
            14'h0879: o_data_a = 16'b0000100001111101;
            14'h087a: o_data_a = 16'b1110110000010000;
            14'h087b: o_data_a = 16'b0000000001011111;
            14'h087c: o_data_a = 16'b1110101010000111;
            14'h087d: o_data_a = 16'b0000000000000000;
            14'h087e: o_data_a = 16'b1111110010101000;
            14'h087f: o_data_a = 16'b1111110000010000;
            14'h0880: o_data_a = 16'b0000000000000001;
            14'h0881: o_data_a = 16'b1111110111100000;
            14'h0882: o_data_a = 16'b1110001100001000;
            14'h0883: o_data_a = 16'b0000000000000011;
            14'h0884: o_data_a = 16'b1111110111100000;
            14'h0885: o_data_a = 16'b1111110000010000;
            14'h0886: o_data_a = 16'b0000000000000000;
            14'h0887: o_data_a = 16'b1111110111101000;
            14'h0888: o_data_a = 16'b1110110010100000;
            14'h0889: o_data_a = 16'b1110001100001000;
            14'h088a: o_data_a = 16'b0000000000000001;
            14'h088b: o_data_a = 16'b1111110111100000;
            14'h088c: o_data_a = 16'b1111110000010000;
            14'h088d: o_data_a = 16'b0000000000000000;
            14'h088e: o_data_a = 16'b1111110111101000;
            14'h088f: o_data_a = 16'b1110110010100000;
            14'h0890: o_data_a = 16'b1110001100001000;
            14'h0891: o_data_a = 16'b0000000000000001;
            14'h0892: o_data_a = 16'b1111110000010000;
            14'h0893: o_data_a = 16'b0000000000000100;
            14'h0894: o_data_a = 16'b1110000010100000;
            14'h0895: o_data_a = 16'b1111110000010000;
            14'h0896: o_data_a = 16'b0000000000000000;
            14'h0897: o_data_a = 16'b1111110111101000;
            14'h0898: o_data_a = 16'b1110110010100000;
            14'h0899: o_data_a = 16'b1110001100001000;
            14'h089a: o_data_a = 16'b0000000000000010;
            14'h089b: o_data_a = 16'b1110110000010000;
            14'h089c: o_data_a = 16'b0000000000001101;
            14'h089d: o_data_a = 16'b1110001100001000;
            14'h089e: o_data_a = 16'b0001101010100110;
            14'h089f: o_data_a = 16'b1110110000010000;
            14'h08a0: o_data_a = 16'b0000000000001110;
            14'h08a1: o_data_a = 16'b1110001100001000;
            14'h08a2: o_data_a = 16'b0000100010100110;
            14'h08a3: o_data_a = 16'b1110110000010000;
            14'h08a4: o_data_a = 16'b0000000001011111;
            14'h08a5: o_data_a = 16'b1110101010000111;
            14'h08a6: o_data_a = 16'b0000000000000000;
            14'h08a7: o_data_a = 16'b1111110010101000;
            14'h08a8: o_data_a = 16'b1111110000010000;
            14'h08a9: o_data_a = 16'b1110110010100000;
            14'h08aa: o_data_a = 16'b1111000010001000;
            14'h08ab: o_data_a = 16'b0000000000000000;
            14'h08ac: o_data_a = 16'b1111110010101000;
            14'h08ad: o_data_a = 16'b1111110000010000;
            14'h08ae: o_data_a = 16'b0000000000000001;
            14'h08af: o_data_a = 16'b1111110111100000;
            14'h08b0: o_data_a = 16'b1110001100001000;
            14'h08b1: o_data_a = 16'b0000101000111000;
            14'h08b2: o_data_a = 16'b1110101010000111;
            14'h08b3: o_data_a = 16'b0000000000000011;
            14'h08b4: o_data_a = 16'b1111110000010000;
            14'h08b5: o_data_a = 16'b0000000000001110;
            14'h08b6: o_data_a = 16'b1110000010100000;
            14'h08b7: o_data_a = 16'b1111110000010000;
            14'h08b8: o_data_a = 16'b0000000000000000;
            14'h08b9: o_data_a = 16'b1111110111101000;
            14'h08ba: o_data_a = 16'b1110110010100000;
            14'h08bb: o_data_a = 16'b1110001100001000;
            14'h08bc: o_data_a = 16'b0000000000000010;
            14'h08bd: o_data_a = 16'b1110110000010000;
            14'h08be: o_data_a = 16'b0000000000000000;
            14'h08bf: o_data_a = 16'b1111110111101000;
            14'h08c0: o_data_a = 16'b1110110010100000;
            14'h08c1: o_data_a = 16'b1110001100001000;
            14'h08c2: o_data_a = 16'b0000100011000110;
            14'h08c3: o_data_a = 16'b1110110000010000;
            14'h08c4: o_data_a = 16'b0000000000000110;
            14'h08c5: o_data_a = 16'b1110101010000111;
            14'h08c6: o_data_a = 16'b0000000000000000;
            14'h08c7: o_data_a = 16'b1111110010101000;
            14'h08c8: o_data_a = 16'b1111110000010000;
            14'h08c9: o_data_a = 16'b0000100011001101;
            14'h08ca: o_data_a = 16'b1110001100000101;
            14'h08cb: o_data_a = 16'b0000100100111100;
            14'h08cc: o_data_a = 16'b1110101010000111;
            14'h08cd: o_data_a = 16'b0000000000000000;
            14'h08ce: o_data_a = 16'b1111110111001000;
            14'h08cf: o_data_a = 16'b1111110010100000;
            14'h08d0: o_data_a = 16'b1110101010001000;
            14'h08d1: o_data_a = 16'b0000000000000000;
            14'h08d2: o_data_a = 16'b1111110010101000;
            14'h08d3: o_data_a = 16'b1111110000010000;
            14'h08d4: o_data_a = 16'b0000000000000001;
            14'h08d5: o_data_a = 16'b1111110000100000;
            14'h08d6: o_data_a = 16'b1110001100001000;
            14'h08d7: o_data_a = 16'b0000000000000001;
            14'h08d8: o_data_a = 16'b1111110000010000;
            14'h08d9: o_data_a = 16'b0000000000000011;
            14'h08da: o_data_a = 16'b1110000010100000;
            14'h08db: o_data_a = 16'b1111110000010000;
            14'h08dc: o_data_a = 16'b0000000000000000;
            14'h08dd: o_data_a = 16'b1111110111101000;
            14'h08de: o_data_a = 16'b1110110010100000;
            14'h08df: o_data_a = 16'b1110001100001000;
            14'h08e0: o_data_a = 16'b0000000000110010;
            14'h08e1: o_data_a = 16'b1110110000010000;
            14'h08e2: o_data_a = 16'b0000000000000000;
            14'h08e3: o_data_a = 16'b1111110111101000;
            14'h08e4: o_data_a = 16'b1110110010100000;
            14'h08e5: o_data_a = 16'b1110001100001000;
            14'h08e6: o_data_a = 16'b0000000000000010;
            14'h08e7: o_data_a = 16'b1110110000010000;
            14'h08e8: o_data_a = 16'b0000000000001101;
            14'h08e9: o_data_a = 16'b1110001100001000;
            14'h08ea: o_data_a = 16'b0001101010100110;
            14'h08eb: o_data_a = 16'b1110110000010000;
            14'h08ec: o_data_a = 16'b0000000000001110;
            14'h08ed: o_data_a = 16'b1110001100001000;
            14'h08ee: o_data_a = 16'b0000100011110010;
            14'h08ef: o_data_a = 16'b1110110000010000;
            14'h08f0: o_data_a = 16'b0000000001011111;
            14'h08f1: o_data_a = 16'b1110101010000111;
            14'h08f2: o_data_a = 16'b0000000000000001;
            14'h08f3: o_data_a = 16'b1111110111100000;
            14'h08f4: o_data_a = 16'b1110110111100000;
            14'h08f5: o_data_a = 16'b1111110000010000;
            14'h08f6: o_data_a = 16'b0000000000000000;
            14'h08f7: o_data_a = 16'b1111110111101000;
            14'h08f8: o_data_a = 16'b1110110010100000;
            14'h08f9: o_data_a = 16'b1110001100001000;
            14'h08fa: o_data_a = 16'b0000000000000010;
            14'h08fb: o_data_a = 16'b1110110000010000;
            14'h08fc: o_data_a = 16'b0000000000001101;
            14'h08fd: o_data_a = 16'b1110001100001000;
            14'h08fe: o_data_a = 16'b0001110001110111;
            14'h08ff: o_data_a = 16'b1110110000010000;
            14'h0900: o_data_a = 16'b0000000000001110;
            14'h0901: o_data_a = 16'b1110001100001000;
            14'h0902: o_data_a = 16'b0000100100000110;
            14'h0903: o_data_a = 16'b1110110000010000;
            14'h0904: o_data_a = 16'b0000000001011111;
            14'h0905: o_data_a = 16'b1110101010000111;
            14'h0906: o_data_a = 16'b0000000000000000;
            14'h0907: o_data_a = 16'b1111110010101000;
            14'h0908: o_data_a = 16'b1111110000010000;
            14'h0909: o_data_a = 16'b0000000000000001;
            14'h090a: o_data_a = 16'b1111110111100000;
            14'h090b: o_data_a = 16'b1110001100001000;
            14'h090c: o_data_a = 16'b0000000000000011;
            14'h090d: o_data_a = 16'b1111110111100000;
            14'h090e: o_data_a = 16'b1111110000010000;
            14'h090f: o_data_a = 16'b0000000000000000;
            14'h0910: o_data_a = 16'b1111110111101000;
            14'h0911: o_data_a = 16'b1110110010100000;
            14'h0912: o_data_a = 16'b1110001100001000;
            14'h0913: o_data_a = 16'b0000000000000001;
            14'h0914: o_data_a = 16'b1111110111100000;
            14'h0915: o_data_a = 16'b1111110000010000;
            14'h0916: o_data_a = 16'b0000000000000000;
            14'h0917: o_data_a = 16'b1111110111101000;
            14'h0918: o_data_a = 16'b1110110010100000;
            14'h0919: o_data_a = 16'b1110001100001000;
            14'h091a: o_data_a = 16'b0000000000000001;
            14'h091b: o_data_a = 16'b1111110000010000;
            14'h091c: o_data_a = 16'b0000000000000100;
            14'h091d: o_data_a = 16'b1110000010100000;
            14'h091e: o_data_a = 16'b1111110000010000;
            14'h091f: o_data_a = 16'b0000000000000000;
            14'h0920: o_data_a = 16'b1111110111101000;
            14'h0921: o_data_a = 16'b1110110010100000;
            14'h0922: o_data_a = 16'b1110001100001000;
            14'h0923: o_data_a = 16'b0000000000000010;
            14'h0924: o_data_a = 16'b1110110000010000;
            14'h0925: o_data_a = 16'b0000000000001101;
            14'h0926: o_data_a = 16'b1110001100001000;
            14'h0927: o_data_a = 16'b0001101010100110;
            14'h0928: o_data_a = 16'b1110110000010000;
            14'h0929: o_data_a = 16'b0000000000001110;
            14'h092a: o_data_a = 16'b1110001100001000;
            14'h092b: o_data_a = 16'b0000100100101111;
            14'h092c: o_data_a = 16'b1110110000010000;
            14'h092d: o_data_a = 16'b0000000001011111;
            14'h092e: o_data_a = 16'b1110101010000111;
            14'h092f: o_data_a = 16'b0000000000000000;
            14'h0930: o_data_a = 16'b1111110010101000;
            14'h0931: o_data_a = 16'b1111110000010000;
            14'h0932: o_data_a = 16'b1110110010100000;
            14'h0933: o_data_a = 16'b1111000010001000;
            14'h0934: o_data_a = 16'b0000000000000000;
            14'h0935: o_data_a = 16'b1111110010101000;
            14'h0936: o_data_a = 16'b1111110000010000;
            14'h0937: o_data_a = 16'b0000000000000001;
            14'h0938: o_data_a = 16'b1111110111100000;
            14'h0939: o_data_a = 16'b1110001100001000;
            14'h093a: o_data_a = 16'b0000101000111000;
            14'h093b: o_data_a = 16'b1110101010000111;
            14'h093c: o_data_a = 16'b0000000000000011;
            14'h093d: o_data_a = 16'b1111110000010000;
            14'h093e: o_data_a = 16'b0000000000001110;
            14'h093f: o_data_a = 16'b1110000010100000;
            14'h0940: o_data_a = 16'b1111110000010000;
            14'h0941: o_data_a = 16'b0000000000000000;
            14'h0942: o_data_a = 16'b1111110111101000;
            14'h0943: o_data_a = 16'b1110110010100000;
            14'h0944: o_data_a = 16'b1110001100001000;
            14'h0945: o_data_a = 16'b0000000000000011;
            14'h0946: o_data_a = 16'b1110110000010000;
            14'h0947: o_data_a = 16'b0000000000000000;
            14'h0948: o_data_a = 16'b1111110111101000;
            14'h0949: o_data_a = 16'b1110110010100000;
            14'h094a: o_data_a = 16'b1110001100001000;
            14'h094b: o_data_a = 16'b0000100101001111;
            14'h094c: o_data_a = 16'b1110110000010000;
            14'h094d: o_data_a = 16'b0000000000000110;
            14'h094e: o_data_a = 16'b1110101010000111;
            14'h094f: o_data_a = 16'b0000000000000000;
            14'h0950: o_data_a = 16'b1111110010101000;
            14'h0951: o_data_a = 16'b1111110000010000;
            14'h0952: o_data_a = 16'b0000100101010110;
            14'h0953: o_data_a = 16'b1110001100000101;
            14'h0954: o_data_a = 16'b0000100111001011;
            14'h0955: o_data_a = 16'b1110101010000111;
            14'h0956: o_data_a = 16'b0000000011111010;
            14'h0957: o_data_a = 16'b1110110000010000;
            14'h0958: o_data_a = 16'b0000000000000000;
            14'h0959: o_data_a = 16'b1111110111101000;
            14'h095a: o_data_a = 16'b1110110010100000;
            14'h095b: o_data_a = 16'b1110001100001000;
            14'h095c: o_data_a = 16'b0000000000000000;
            14'h095d: o_data_a = 16'b1111110010101000;
            14'h095e: o_data_a = 16'b1111110000010000;
            14'h095f: o_data_a = 16'b0000000000000001;
            14'h0960: o_data_a = 16'b1111110111100000;
            14'h0961: o_data_a = 16'b1110001100001000;
            14'h0962: o_data_a = 16'b0000000000000001;
            14'h0963: o_data_a = 16'b1111110111100000;
            14'h0964: o_data_a = 16'b1110110111100000;
            14'h0965: o_data_a = 16'b1111110000010000;
            14'h0966: o_data_a = 16'b0000000000000000;
            14'h0967: o_data_a = 16'b1111110111101000;
            14'h0968: o_data_a = 16'b1110110010100000;
            14'h0969: o_data_a = 16'b1110001100001000;
            14'h096a: o_data_a = 16'b0000000000011001;
            14'h096b: o_data_a = 16'b1110110000010000;
            14'h096c: o_data_a = 16'b0000000000000000;
            14'h096d: o_data_a = 16'b1111110111101000;
            14'h096e: o_data_a = 16'b1110110010100000;
            14'h096f: o_data_a = 16'b1110001100001000;
            14'h0970: o_data_a = 16'b0000000000000000;
            14'h0971: o_data_a = 16'b1111110010100000;
            14'h0972: o_data_a = 16'b1111110001010000;
            14'h0973: o_data_a = 16'b1110011111001000;
            14'h0974: o_data_a = 16'b0000000000000010;
            14'h0975: o_data_a = 16'b1110110000010000;
            14'h0976: o_data_a = 16'b0000000000001101;
            14'h0977: o_data_a = 16'b1110001100001000;
            14'h0978: o_data_a = 16'b0001101010100110;
            14'h0979: o_data_a = 16'b1110110000010000;
            14'h097a: o_data_a = 16'b0000000000001110;
            14'h097b: o_data_a = 16'b1110001100001000;
            14'h097c: o_data_a = 16'b0000100110000000;
            14'h097d: o_data_a = 16'b1110110000010000;
            14'h097e: o_data_a = 16'b0000000001011111;
            14'h097f: o_data_a = 16'b1110101010000111;
            14'h0980: o_data_a = 16'b0000000000000001;
            14'h0981: o_data_a = 16'b1111110000010000;
            14'h0982: o_data_a = 16'b0000000000000011;
            14'h0983: o_data_a = 16'b1110000010100000;
            14'h0984: o_data_a = 16'b1111110000010000;
            14'h0985: o_data_a = 16'b0000000000000000;
            14'h0986: o_data_a = 16'b1111110111101000;
            14'h0987: o_data_a = 16'b1110110010100000;
            14'h0988: o_data_a = 16'b1110001100001000;
            14'h0989: o_data_a = 16'b0000000000000010;
            14'h098a: o_data_a = 16'b1110110000010000;
            14'h098b: o_data_a = 16'b0000000000001101;
            14'h098c: o_data_a = 16'b1110001100001000;
            14'h098d: o_data_a = 16'b0001110001110111;
            14'h098e: o_data_a = 16'b1110110000010000;
            14'h098f: o_data_a = 16'b0000000000001110;
            14'h0990: o_data_a = 16'b1110001100001000;
            14'h0991: o_data_a = 16'b0000100110010101;
            14'h0992: o_data_a = 16'b1110110000010000;
            14'h0993: o_data_a = 16'b0000000001011111;
            14'h0994: o_data_a = 16'b1110101010000111;
            14'h0995: o_data_a = 16'b0000000000000000;
            14'h0996: o_data_a = 16'b1111110010101000;
            14'h0997: o_data_a = 16'b1111110000010000;
            14'h0998: o_data_a = 16'b0000000000000001;
            14'h0999: o_data_a = 16'b1111110000100000;
            14'h099a: o_data_a = 16'b1110001100001000;
            14'h099b: o_data_a = 16'b0000000000000011;
            14'h099c: o_data_a = 16'b1111110000100000;
            14'h099d: o_data_a = 16'b1111110000010000;
            14'h099e: o_data_a = 16'b0000000000000000;
            14'h099f: o_data_a = 16'b1111110111101000;
            14'h09a0: o_data_a = 16'b1110110010100000;
            14'h09a1: o_data_a = 16'b1110001100001000;
            14'h09a2: o_data_a = 16'b0000000000000001;
            14'h09a3: o_data_a = 16'b1111110000100000;
            14'h09a4: o_data_a = 16'b1111110000010000;
            14'h09a5: o_data_a = 16'b0000000000000000;
            14'h09a6: o_data_a = 16'b1111110111101000;
            14'h09a7: o_data_a = 16'b1110110010100000;
            14'h09a8: o_data_a = 16'b1110001100001000;
            14'h09a9: o_data_a = 16'b0000000000000001;
            14'h09aa: o_data_a = 16'b1111110000010000;
            14'h09ab: o_data_a = 16'b0000000000000100;
            14'h09ac: o_data_a = 16'b1110000010100000;
            14'h09ad: o_data_a = 16'b1111110000010000;
            14'h09ae: o_data_a = 16'b0000000000000000;
            14'h09af: o_data_a = 16'b1111110111101000;
            14'h09b0: o_data_a = 16'b1110110010100000;
            14'h09b1: o_data_a = 16'b1110001100001000;
            14'h09b2: o_data_a = 16'b0000000000000010;
            14'h09b3: o_data_a = 16'b1110110000010000;
            14'h09b4: o_data_a = 16'b0000000000001101;
            14'h09b5: o_data_a = 16'b1110001100001000;
            14'h09b6: o_data_a = 16'b0001101010100110;
            14'h09b7: o_data_a = 16'b1110110000010000;
            14'h09b8: o_data_a = 16'b0000000000001110;
            14'h09b9: o_data_a = 16'b1110001100001000;
            14'h09ba: o_data_a = 16'b0000100110111110;
            14'h09bb: o_data_a = 16'b1110110000010000;
            14'h09bc: o_data_a = 16'b0000000001011111;
            14'h09bd: o_data_a = 16'b1110101010000111;
            14'h09be: o_data_a = 16'b0000000000000000;
            14'h09bf: o_data_a = 16'b1111110010101000;
            14'h09c0: o_data_a = 16'b1111110000010000;
            14'h09c1: o_data_a = 16'b1110110010100000;
            14'h09c2: o_data_a = 16'b1111000010001000;
            14'h09c3: o_data_a = 16'b0000000000000000;
            14'h09c4: o_data_a = 16'b1111110010101000;
            14'h09c5: o_data_a = 16'b1111110000010000;
            14'h09c6: o_data_a = 16'b0000000000000001;
            14'h09c7: o_data_a = 16'b1111110000100000;
            14'h09c8: o_data_a = 16'b1110001100001000;
            14'h09c9: o_data_a = 16'b0000101000111000;
            14'h09ca: o_data_a = 16'b1110101010000111;
            14'h09cb: o_data_a = 16'b0000000000000000;
            14'h09cc: o_data_a = 16'b1111110111001000;
            14'h09cd: o_data_a = 16'b1111110010100000;
            14'h09ce: o_data_a = 16'b1110101010001000;
            14'h09cf: o_data_a = 16'b0000000000000000;
            14'h09d0: o_data_a = 16'b1111110010101000;
            14'h09d1: o_data_a = 16'b1111110000010000;
            14'h09d2: o_data_a = 16'b0000000000000001;
            14'h09d3: o_data_a = 16'b1111110111100000;
            14'h09d4: o_data_a = 16'b1110001100001000;
            14'h09d5: o_data_a = 16'b0000000000000001;
            14'h09d6: o_data_a = 16'b1111110111100000;
            14'h09d7: o_data_a = 16'b1110110111100000;
            14'h09d8: o_data_a = 16'b1111110000010000;
            14'h09d9: o_data_a = 16'b0000000000000000;
            14'h09da: o_data_a = 16'b1111110111101000;
            14'h09db: o_data_a = 16'b1110110010100000;
            14'h09dc: o_data_a = 16'b1110001100001000;
            14'h09dd: o_data_a = 16'b0000000000011001;
            14'h09de: o_data_a = 16'b1110110000010000;
            14'h09df: o_data_a = 16'b0000000000000000;
            14'h09e0: o_data_a = 16'b1111110111101000;
            14'h09e1: o_data_a = 16'b1110110010100000;
            14'h09e2: o_data_a = 16'b1110001100001000;
            14'h09e3: o_data_a = 16'b0000000000000010;
            14'h09e4: o_data_a = 16'b1110110000010000;
            14'h09e5: o_data_a = 16'b0000000000001101;
            14'h09e6: o_data_a = 16'b1110001100001000;
            14'h09e7: o_data_a = 16'b0001101010100110;
            14'h09e8: o_data_a = 16'b1110110000010000;
            14'h09e9: o_data_a = 16'b0000000000001110;
            14'h09ea: o_data_a = 16'b1110001100001000;
            14'h09eb: o_data_a = 16'b0000100111101111;
            14'h09ec: o_data_a = 16'b1110110000010000;
            14'h09ed: o_data_a = 16'b0000000001011111;
            14'h09ee: o_data_a = 16'b1110101010000111;
            14'h09ef: o_data_a = 16'b0000000000000001;
            14'h09f0: o_data_a = 16'b1111110000010000;
            14'h09f1: o_data_a = 16'b0000000000000011;
            14'h09f2: o_data_a = 16'b1110000010100000;
            14'h09f3: o_data_a = 16'b1111110000010000;
            14'h09f4: o_data_a = 16'b0000000000000000;
            14'h09f5: o_data_a = 16'b1111110111101000;
            14'h09f6: o_data_a = 16'b1110110010100000;
            14'h09f7: o_data_a = 16'b1110001100001000;
            14'h09f8: o_data_a = 16'b0000000000000010;
            14'h09f9: o_data_a = 16'b1110110000010000;
            14'h09fa: o_data_a = 16'b0000000000001101;
            14'h09fb: o_data_a = 16'b1110001100001000;
            14'h09fc: o_data_a = 16'b0001110001110111;
            14'h09fd: o_data_a = 16'b1110110000010000;
            14'h09fe: o_data_a = 16'b0000000000001110;
            14'h09ff: o_data_a = 16'b1110001100001000;
            14'h0a00: o_data_a = 16'b0000101000000100;
            14'h0a01: o_data_a = 16'b1110110000010000;
            14'h0a02: o_data_a = 16'b0000000001011111;
            14'h0a03: o_data_a = 16'b1110101010000111;
            14'h0a04: o_data_a = 16'b0000000000000000;
            14'h0a05: o_data_a = 16'b1111110010101000;
            14'h0a06: o_data_a = 16'b1111110000010000;
            14'h0a07: o_data_a = 16'b0000000000000001;
            14'h0a08: o_data_a = 16'b1111110000100000;
            14'h0a09: o_data_a = 16'b1110001100001000;
            14'h0a0a: o_data_a = 16'b0000000000000011;
            14'h0a0b: o_data_a = 16'b1111110000100000;
            14'h0a0c: o_data_a = 16'b1111110000010000;
            14'h0a0d: o_data_a = 16'b0000000000000000;
            14'h0a0e: o_data_a = 16'b1111110111101000;
            14'h0a0f: o_data_a = 16'b1110110010100000;
            14'h0a10: o_data_a = 16'b1110001100001000;
            14'h0a11: o_data_a = 16'b0000000000000001;
            14'h0a12: o_data_a = 16'b1111110000100000;
            14'h0a13: o_data_a = 16'b1111110000010000;
            14'h0a14: o_data_a = 16'b0000000000000000;
            14'h0a15: o_data_a = 16'b1111110111101000;
            14'h0a16: o_data_a = 16'b1110110010100000;
            14'h0a17: o_data_a = 16'b1110001100001000;
            14'h0a18: o_data_a = 16'b0000000000000001;
            14'h0a19: o_data_a = 16'b1111110000010000;
            14'h0a1a: o_data_a = 16'b0000000000000100;
            14'h0a1b: o_data_a = 16'b1110000010100000;
            14'h0a1c: o_data_a = 16'b1111110000010000;
            14'h0a1d: o_data_a = 16'b0000000000000000;
            14'h0a1e: o_data_a = 16'b1111110111101000;
            14'h0a1f: o_data_a = 16'b1110110010100000;
            14'h0a20: o_data_a = 16'b1110001100001000;
            14'h0a21: o_data_a = 16'b0000000000000010;
            14'h0a22: o_data_a = 16'b1110110000010000;
            14'h0a23: o_data_a = 16'b0000000000001101;
            14'h0a24: o_data_a = 16'b1110001100001000;
            14'h0a25: o_data_a = 16'b0001101010100110;
            14'h0a26: o_data_a = 16'b1110110000010000;
            14'h0a27: o_data_a = 16'b0000000000001110;
            14'h0a28: o_data_a = 16'b1110001100001000;
            14'h0a29: o_data_a = 16'b0000101000101101;
            14'h0a2a: o_data_a = 16'b1110110000010000;
            14'h0a2b: o_data_a = 16'b0000000001011111;
            14'h0a2c: o_data_a = 16'b1110101010000111;
            14'h0a2d: o_data_a = 16'b0000000000000000;
            14'h0a2e: o_data_a = 16'b1111110010101000;
            14'h0a2f: o_data_a = 16'b1111110000010000;
            14'h0a30: o_data_a = 16'b1110110010100000;
            14'h0a31: o_data_a = 16'b1111000010001000;
            14'h0a32: o_data_a = 16'b0000000000000000;
            14'h0a33: o_data_a = 16'b1111110010101000;
            14'h0a34: o_data_a = 16'b1111110000010000;
            14'h0a35: o_data_a = 16'b0000000000000001;
            14'h0a36: o_data_a = 16'b1111110000100000;
            14'h0a37: o_data_a = 16'b1110001100001000;
            14'h0a38: o_data_a = 16'b0000000000000011;
            14'h0a39: o_data_a = 16'b1111110000010000;
            14'h0a3a: o_data_a = 16'b0000000000000000;
            14'h0a3b: o_data_a = 16'b1111110111101000;
            14'h0a3c: o_data_a = 16'b1110110010100000;
            14'h0a3d: o_data_a = 16'b1110001100001000;
            14'h0a3e: o_data_a = 16'b0000000000000001;
            14'h0a3f: o_data_a = 16'b1111110000100000;
            14'h0a40: o_data_a = 16'b1111110000010000;
            14'h0a41: o_data_a = 16'b0000000000000000;
            14'h0a42: o_data_a = 16'b1111110111101000;
            14'h0a43: o_data_a = 16'b1110110010100000;
            14'h0a44: o_data_a = 16'b1110001100001000;
            14'h0a45: o_data_a = 16'b0000000000000001;
            14'h0a46: o_data_a = 16'b1111110111100000;
            14'h0a47: o_data_a = 16'b1111110000010000;
            14'h0a48: o_data_a = 16'b0000000000000000;
            14'h0a49: o_data_a = 16'b1111110111101000;
            14'h0a4a: o_data_a = 16'b1110110010100000;
            14'h0a4b: o_data_a = 16'b1110001100001000;
            14'h0a4c: o_data_a = 16'b0000000000000011;
            14'h0a4d: o_data_a = 16'b1110110000010000;
            14'h0a4e: o_data_a = 16'b0000000000001101;
            14'h0a4f: o_data_a = 16'b1110001100001000;
            14'h0a50: o_data_a = 16'b0000001010001100;
            14'h0a51: o_data_a = 16'b1110110000010000;
            14'h0a52: o_data_a = 16'b0000000000001110;
            14'h0a53: o_data_a = 16'b1110001100001000;
            14'h0a54: o_data_a = 16'b0000101001011000;
            14'h0a55: o_data_a = 16'b1110110000010000;
            14'h0a56: o_data_a = 16'b0000000001011111;
            14'h0a57: o_data_a = 16'b1110101010000111;
            14'h0a58: o_data_a = 16'b0000000000000000;
            14'h0a59: o_data_a = 16'b1111110010101000;
            14'h0a5a: o_data_a = 16'b1111110000010000;
            14'h0a5b: o_data_a = 16'b0000000000000101;
            14'h0a5c: o_data_a = 16'b1110001100001000;
            14'h0a5d: o_data_a = 16'b0000000000000000;
            14'h0a5e: o_data_a = 16'b1111110111001000;
            14'h0a5f: o_data_a = 16'b1111110010100000;
            14'h0a60: o_data_a = 16'b1110101010001000;
            14'h0a61: o_data_a = 16'b0000000000110110;
            14'h0a62: o_data_a = 16'b1110101010000111;
            14'h0a63: o_data_a = 16'b0000000000000101;
            14'h0a64: o_data_a = 16'b1110110000010000;
            14'h0a65: o_data_a = 16'b0000000000000000;
            14'h0a66: o_data_a = 16'b1111110111101000;
            14'h0a67: o_data_a = 16'b1110110010100000;
            14'h0a68: o_data_a = 16'b1110001100001000;
            14'h0a69: o_data_a = 16'b0000000000000001;
            14'h0a6a: o_data_a = 16'b1110110000010000;
            14'h0a6b: o_data_a = 16'b0000000000001101;
            14'h0a6c: o_data_a = 16'b1110001100001000;
            14'h0a6d: o_data_a = 16'b0010000111000011;
            14'h0a6e: o_data_a = 16'b1110110000010000;
            14'h0a6f: o_data_a = 16'b0000000000001110;
            14'h0a70: o_data_a = 16'b1110001100001000;
            14'h0a71: o_data_a = 16'b0000101001110101;
            14'h0a72: o_data_a = 16'b1110110000010000;
            14'h0a73: o_data_a = 16'b0000000001011111;
            14'h0a74: o_data_a = 16'b1110101010000111;
            14'h0a75: o_data_a = 16'b0000000000000000;
            14'h0a76: o_data_a = 16'b1111110010101000;
            14'h0a77: o_data_a = 16'b1111110000010000;
            14'h0a78: o_data_a = 16'b0000000000000011;
            14'h0a79: o_data_a = 16'b1110001100001000;
            14'h0a7a: o_data_a = 16'b0000000000000010;
            14'h0a7b: o_data_a = 16'b1111110000100000;
            14'h0a7c: o_data_a = 16'b1111110000010000;
            14'h0a7d: o_data_a = 16'b0000000000000000;
            14'h0a7e: o_data_a = 16'b1111110111101000;
            14'h0a7f: o_data_a = 16'b1110110010100000;
            14'h0a80: o_data_a = 16'b1110001100001000;
            14'h0a81: o_data_a = 16'b0000000000000000;
            14'h0a82: o_data_a = 16'b1111110010101000;
            14'h0a83: o_data_a = 16'b1111110000010000;
            14'h0a84: o_data_a = 16'b0000000000000011;
            14'h0a85: o_data_a = 16'b1111110000100000;
            14'h0a86: o_data_a = 16'b1110001100001000;
            14'h0a87: o_data_a = 16'b0000000000000010;
            14'h0a88: o_data_a = 16'b1111110111100000;
            14'h0a89: o_data_a = 16'b1111110000010000;
            14'h0a8a: o_data_a = 16'b0000000000000000;
            14'h0a8b: o_data_a = 16'b1111110111101000;
            14'h0a8c: o_data_a = 16'b1110110010100000;
            14'h0a8d: o_data_a = 16'b1110001100001000;
            14'h0a8e: o_data_a = 16'b0000000000000000;
            14'h0a8f: o_data_a = 16'b1111110010101000;
            14'h0a90: o_data_a = 16'b1111110000010000;
            14'h0a91: o_data_a = 16'b0000000000000011;
            14'h0a92: o_data_a = 16'b1111110111100000;
            14'h0a93: o_data_a = 16'b1110001100001000;
            14'h0a94: o_data_a = 16'b0000000000000010;
            14'h0a95: o_data_a = 16'b1111110111100000;
            14'h0a96: o_data_a = 16'b1110110111100000;
            14'h0a97: o_data_a = 16'b1111110000010000;
            14'h0a98: o_data_a = 16'b0000000000000000;
            14'h0a99: o_data_a = 16'b1111110111101000;
            14'h0a9a: o_data_a = 16'b1110110010100000;
            14'h0a9b: o_data_a = 16'b1110001100001000;
            14'h0a9c: o_data_a = 16'b0000000000000000;
            14'h0a9d: o_data_a = 16'b1111110010101000;
            14'h0a9e: o_data_a = 16'b1111110000010000;
            14'h0a9f: o_data_a = 16'b0000000000000011;
            14'h0aa0: o_data_a = 16'b1111110111100000;
            14'h0aa1: o_data_a = 16'b1110110111100000;
            14'h0aa2: o_data_a = 16'b1110001100001000;
            14'h0aa3: o_data_a = 16'b0000000000000010;
            14'h0aa4: o_data_a = 16'b1111110000010000;
            14'h0aa5: o_data_a = 16'b0000000000000011;
            14'h0aa6: o_data_a = 16'b1110000010100000;
            14'h0aa7: o_data_a = 16'b1111110000010000;
            14'h0aa8: o_data_a = 16'b0000000000000000;
            14'h0aa9: o_data_a = 16'b1111110111101000;
            14'h0aaa: o_data_a = 16'b1110110010100000;
            14'h0aab: o_data_a = 16'b1110001100001000;
            14'h0aac: o_data_a = 16'b0000000000000000;
            14'h0aad: o_data_a = 16'b1111110010101000;
            14'h0aae: o_data_a = 16'b1111110000010000;
            14'h0aaf: o_data_a = 16'b0000000000000011;
            14'h0ab0: o_data_a = 16'b1111110111100000;
            14'h0ab1: o_data_a = 16'b1110110111100000;
            14'h0ab2: o_data_a = 16'b1110110111100000;
            14'h0ab3: o_data_a = 16'b1110001100001000;
            14'h0ab4: o_data_a = 16'b0000000000000010;
            14'h0ab5: o_data_a = 16'b1110110000010000;
            14'h0ab6: o_data_a = 16'b0000000000000000;
            14'h0ab7: o_data_a = 16'b1111110111101000;
            14'h0ab8: o_data_a = 16'b1110110010100000;
            14'h0ab9: o_data_a = 16'b1110001100001000;
            14'h0aba: o_data_a = 16'b0000000000000000;
            14'h0abb: o_data_a = 16'b1111110010101000;
            14'h0abc: o_data_a = 16'b1111110000010000;
            14'h0abd: o_data_a = 16'b0000000000000011;
            14'h0abe: o_data_a = 16'b1111110111100000;
            14'h0abf: o_data_a = 16'b1110110111100000;
            14'h0ac0: o_data_a = 16'b1110110111100000;
            14'h0ac1: o_data_a = 16'b1110110111100000;
            14'h0ac2: o_data_a = 16'b1110001100001000;
            14'h0ac3: o_data_a = 16'b0000000000000011;
            14'h0ac4: o_data_a = 16'b1111110000010000;
            14'h0ac5: o_data_a = 16'b0000000000000000;
            14'h0ac6: o_data_a = 16'b1111110111101000;
            14'h0ac7: o_data_a = 16'b1110110010100000;
            14'h0ac8: o_data_a = 16'b1110001100001000;
            14'h0ac9: o_data_a = 16'b0000000000000001;
            14'h0aca: o_data_a = 16'b1110110000010000;
            14'h0acb: o_data_a = 16'b0000000000001101;
            14'h0acc: o_data_a = 16'b1110001100001000;
            14'h0acd: o_data_a = 16'b0000101100001011;
            14'h0ace: o_data_a = 16'b1110110000010000;
            14'h0acf: o_data_a = 16'b0000000000001110;
            14'h0ad0: o_data_a = 16'b1110001100001000;
            14'h0ad1: o_data_a = 16'b0000101011010101;
            14'h0ad2: o_data_a = 16'b1110110000010000;
            14'h0ad3: o_data_a = 16'b0000000001011111;
            14'h0ad4: o_data_a = 16'b1110101010000111;
            14'h0ad5: o_data_a = 16'b0000000000000000;
            14'h0ad6: o_data_a = 16'b1111110010101000;
            14'h0ad7: o_data_a = 16'b1111110000010000;
            14'h0ad8: o_data_a = 16'b0000000000000101;
            14'h0ad9: o_data_a = 16'b1110001100001000;
            14'h0ada: o_data_a = 16'b0000000000000011;
            14'h0adb: o_data_a = 16'b1111110000010000;
            14'h0adc: o_data_a = 16'b0000000000000000;
            14'h0add: o_data_a = 16'b1111110111101000;
            14'h0ade: o_data_a = 16'b1110110010100000;
            14'h0adf: o_data_a = 16'b1110001100001000;
            14'h0ae0: o_data_a = 16'b0000000000110110;
            14'h0ae1: o_data_a = 16'b1110101010000111;
            14'h0ae2: o_data_a = 16'b0000000000000010;
            14'h0ae3: o_data_a = 16'b1111110000100000;
            14'h0ae4: o_data_a = 16'b1111110000010000;
            14'h0ae5: o_data_a = 16'b0000000000000000;
            14'h0ae6: o_data_a = 16'b1111110111101000;
            14'h0ae7: o_data_a = 16'b1110110010100000;
            14'h0ae8: o_data_a = 16'b1110001100001000;
            14'h0ae9: o_data_a = 16'b0000000000000000;
            14'h0aea: o_data_a = 16'b1111110010101000;
            14'h0aeb: o_data_a = 16'b1111110000010000;
            14'h0aec: o_data_a = 16'b0000000000000011;
            14'h0aed: o_data_a = 16'b1110001100001000;
            14'h0aee: o_data_a = 16'b0000000000000011;
            14'h0aef: o_data_a = 16'b1111110000010000;
            14'h0af0: o_data_a = 16'b0000000000000000;
            14'h0af1: o_data_a = 16'b1111110111101000;
            14'h0af2: o_data_a = 16'b1110110010100000;
            14'h0af3: o_data_a = 16'b1110001100001000;
            14'h0af4: o_data_a = 16'b0000000000000001;
            14'h0af5: o_data_a = 16'b1110110000010000;
            14'h0af6: o_data_a = 16'b0000000000001101;
            14'h0af7: o_data_a = 16'b1110001100001000;
            14'h0af8: o_data_a = 16'b0010010010001101;
            14'h0af9: o_data_a = 16'b1110110000010000;
            14'h0afa: o_data_a = 16'b0000000000001110;
            14'h0afb: o_data_a = 16'b1110001100001000;
            14'h0afc: o_data_a = 16'b0000101100000000;
            14'h0afd: o_data_a = 16'b1110110000010000;
            14'h0afe: o_data_a = 16'b0000000001011111;
            14'h0aff: o_data_a = 16'b1110101010000111;
            14'h0b00: o_data_a = 16'b0000000000000000;
            14'h0b01: o_data_a = 16'b1111110010101000;
            14'h0b02: o_data_a = 16'b1111110000010000;
            14'h0b03: o_data_a = 16'b0000000000000101;
            14'h0b04: o_data_a = 16'b1110001100001000;
            14'h0b05: o_data_a = 16'b0000000000000000;
            14'h0b06: o_data_a = 16'b1111110111001000;
            14'h0b07: o_data_a = 16'b1111110010100000;
            14'h0b08: o_data_a = 16'b1110101010001000;
            14'h0b09: o_data_a = 16'b0000000000110110;
            14'h0b0a: o_data_a = 16'b1110101010000111;
            14'h0b0b: o_data_a = 16'b0000000000000010;
            14'h0b0c: o_data_a = 16'b1111110000100000;
            14'h0b0d: o_data_a = 16'b1111110000010000;
            14'h0b0e: o_data_a = 16'b0000000000000000;
            14'h0b0f: o_data_a = 16'b1111110111101000;
            14'h0b10: o_data_a = 16'b1110110010100000;
            14'h0b11: o_data_a = 16'b1110001100001000;
            14'h0b12: o_data_a = 16'b0000000000000000;
            14'h0b13: o_data_a = 16'b1111110010101000;
            14'h0b14: o_data_a = 16'b1111110000010000;
            14'h0b15: o_data_a = 16'b0000000000000011;
            14'h0b16: o_data_a = 16'b1110001100001000;
            14'h0b17: o_data_a = 16'b0000000000000000;
            14'h0b18: o_data_a = 16'b1111110111001000;
            14'h0b19: o_data_a = 16'b1111110010100000;
            14'h0b1a: o_data_a = 16'b1110101010001000;
            14'h0b1b: o_data_a = 16'b0000000000000000;
            14'h0b1c: o_data_a = 16'b1111110010100000;
            14'h0b1d: o_data_a = 16'b1111110001001000;
            14'h0b1e: o_data_a = 16'b0000000000000001;
            14'h0b1f: o_data_a = 16'b1110110000010000;
            14'h0b20: o_data_a = 16'b0000000000001101;
            14'h0b21: o_data_a = 16'b1110001100001000;
            14'h0b22: o_data_a = 16'b0101000110011001;
            14'h0b23: o_data_a = 16'b1110110000010000;
            14'h0b24: o_data_a = 16'b0000000000001110;
            14'h0b25: o_data_a = 16'b1110001100001000;
            14'h0b26: o_data_a = 16'b0000101100101010;
            14'h0b27: o_data_a = 16'b1110110000010000;
            14'h0b28: o_data_a = 16'b0000000001011111;
            14'h0b29: o_data_a = 16'b1110101010000111;
            14'h0b2a: o_data_a = 16'b0000000000000000;
            14'h0b2b: o_data_a = 16'b1111110010101000;
            14'h0b2c: o_data_a = 16'b1111110000010000;
            14'h0b2d: o_data_a = 16'b0000000000000101;
            14'h0b2e: o_data_a = 16'b1110001100001000;
            14'h0b2f: o_data_a = 16'b0000000000000011;
            14'h0b30: o_data_a = 16'b1111110000010000;
            14'h0b31: o_data_a = 16'b0000000000000000;
            14'h0b32: o_data_a = 16'b1111110111101000;
            14'h0b33: o_data_a = 16'b1110110010100000;
            14'h0b34: o_data_a = 16'b1110001100001000;
            14'h0b35: o_data_a = 16'b0000000000000001;
            14'h0b36: o_data_a = 16'b1110110000010000;
            14'h0b37: o_data_a = 16'b0000000000001101;
            14'h0b38: o_data_a = 16'b1110001100001000;
            14'h0b39: o_data_a = 16'b0000101110001010;
            14'h0b3a: o_data_a = 16'b1110110000010000;
            14'h0b3b: o_data_a = 16'b0000000000001110;
            14'h0b3c: o_data_a = 16'b1110001100001000;
            14'h0b3d: o_data_a = 16'b0000101101000001;
            14'h0b3e: o_data_a = 16'b1110110000010000;
            14'h0b3f: o_data_a = 16'b0000000001011111;
            14'h0b40: o_data_a = 16'b1110101010000111;
            14'h0b41: o_data_a = 16'b0000000000000000;
            14'h0b42: o_data_a = 16'b1111110010101000;
            14'h0b43: o_data_a = 16'b1111110000010000;
            14'h0b44: o_data_a = 16'b0000000000000101;
            14'h0b45: o_data_a = 16'b1110001100001000;
            14'h0b46: o_data_a = 16'b0000000000000000;
            14'h0b47: o_data_a = 16'b1111110111001000;
            14'h0b48: o_data_a = 16'b1111110010100000;
            14'h0b49: o_data_a = 16'b1110101010001000;
            14'h0b4a: o_data_a = 16'b0000000000110110;
            14'h0b4b: o_data_a = 16'b1110101010000111;
            14'h0b4c: o_data_a = 16'b0000000000000010;
            14'h0b4d: o_data_a = 16'b1111110000100000;
            14'h0b4e: o_data_a = 16'b1111110000010000;
            14'h0b4f: o_data_a = 16'b0000000000000000;
            14'h0b50: o_data_a = 16'b1111110111101000;
            14'h0b51: o_data_a = 16'b1110110010100000;
            14'h0b52: o_data_a = 16'b1110001100001000;
            14'h0b53: o_data_a = 16'b0000000000000000;
            14'h0b54: o_data_a = 16'b1111110010101000;
            14'h0b55: o_data_a = 16'b1111110000010000;
            14'h0b56: o_data_a = 16'b0000000000000011;
            14'h0b57: o_data_a = 16'b1110001100001000;
            14'h0b58: o_data_a = 16'b0000000000000000;
            14'h0b59: o_data_a = 16'b1111110111001000;
            14'h0b5a: o_data_a = 16'b1111110010100000;
            14'h0b5b: o_data_a = 16'b1110101010001000;
            14'h0b5c: o_data_a = 16'b0000000000000001;
            14'h0b5d: o_data_a = 16'b1110110000010000;
            14'h0b5e: o_data_a = 16'b0000000000001101;
            14'h0b5f: o_data_a = 16'b1110001100001000;
            14'h0b60: o_data_a = 16'b0101000110011001;
            14'h0b61: o_data_a = 16'b1110110000010000;
            14'h0b62: o_data_a = 16'b0000000000001110;
            14'h0b63: o_data_a = 16'b1110001100001000;
            14'h0b64: o_data_a = 16'b0000101101101000;
            14'h0b65: o_data_a = 16'b1110110000010000;
            14'h0b66: o_data_a = 16'b0000000001011111;
            14'h0b67: o_data_a = 16'b1110101010000111;
            14'h0b68: o_data_a = 16'b0000000000000000;
            14'h0b69: o_data_a = 16'b1111110010101000;
            14'h0b6a: o_data_a = 16'b1111110000010000;
            14'h0b6b: o_data_a = 16'b0000000000000101;
            14'h0b6c: o_data_a = 16'b1110001100001000;
            14'h0b6d: o_data_a = 16'b0000000000000011;
            14'h0b6e: o_data_a = 16'b1111110000010000;
            14'h0b6f: o_data_a = 16'b0000000000000000;
            14'h0b70: o_data_a = 16'b1111110111101000;
            14'h0b71: o_data_a = 16'b1110110010100000;
            14'h0b72: o_data_a = 16'b1110001100001000;
            14'h0b73: o_data_a = 16'b0000000000000001;
            14'h0b74: o_data_a = 16'b1110110000010000;
            14'h0b75: o_data_a = 16'b0000000000001101;
            14'h0b76: o_data_a = 16'b1110001100001000;
            14'h0b77: o_data_a = 16'b0000101110001010;
            14'h0b78: o_data_a = 16'b1110110000010000;
            14'h0b79: o_data_a = 16'b0000000000001110;
            14'h0b7a: o_data_a = 16'b1110001100001000;
            14'h0b7b: o_data_a = 16'b0000101101111111;
            14'h0b7c: o_data_a = 16'b1110110000010000;
            14'h0b7d: o_data_a = 16'b0000000001011111;
            14'h0b7e: o_data_a = 16'b1110101010000111;
            14'h0b7f: o_data_a = 16'b0000000000000000;
            14'h0b80: o_data_a = 16'b1111110010101000;
            14'h0b81: o_data_a = 16'b1111110000010000;
            14'h0b82: o_data_a = 16'b0000000000000101;
            14'h0b83: o_data_a = 16'b1110001100001000;
            14'h0b84: o_data_a = 16'b0000000000000000;
            14'h0b85: o_data_a = 16'b1111110111001000;
            14'h0b86: o_data_a = 16'b1111110010100000;
            14'h0b87: o_data_a = 16'b1110101010001000;
            14'h0b88: o_data_a = 16'b0000000000110110;
            14'h0b89: o_data_a = 16'b1110101010000111;
            14'h0b8a: o_data_a = 16'b0000000000000010;
            14'h0b8b: o_data_a = 16'b1111110000100000;
            14'h0b8c: o_data_a = 16'b1111110000010000;
            14'h0b8d: o_data_a = 16'b0000000000000000;
            14'h0b8e: o_data_a = 16'b1111110111101000;
            14'h0b8f: o_data_a = 16'b1110110010100000;
            14'h0b90: o_data_a = 16'b1110001100001000;
            14'h0b91: o_data_a = 16'b0000000000000000;
            14'h0b92: o_data_a = 16'b1111110010101000;
            14'h0b93: o_data_a = 16'b1111110000010000;
            14'h0b94: o_data_a = 16'b0000000000000011;
            14'h0b95: o_data_a = 16'b1110001100001000;
            14'h0b96: o_data_a = 16'b0000000000000011;
            14'h0b97: o_data_a = 16'b1111110000100000;
            14'h0b98: o_data_a = 16'b1111110000010000;
            14'h0b99: o_data_a = 16'b0000000000000000;
            14'h0b9a: o_data_a = 16'b1111110111101000;
            14'h0b9b: o_data_a = 16'b1110110010100000;
            14'h0b9c: o_data_a = 16'b1110001100001000;
            14'h0b9d: o_data_a = 16'b0000000000000011;
            14'h0b9e: o_data_a = 16'b1111110111100000;
            14'h0b9f: o_data_a = 16'b1111110000010000;
            14'h0ba0: o_data_a = 16'b0000000000000000;
            14'h0ba1: o_data_a = 16'b1111110111101000;
            14'h0ba2: o_data_a = 16'b1110110010100000;
            14'h0ba3: o_data_a = 16'b1110001100001000;
            14'h0ba4: o_data_a = 16'b0000000000000011;
            14'h0ba5: o_data_a = 16'b1111110000100000;
            14'h0ba6: o_data_a = 16'b1111110000010000;
            14'h0ba7: o_data_a = 16'b0000000000000000;
            14'h0ba8: o_data_a = 16'b1111110111101000;
            14'h0ba9: o_data_a = 16'b1110110010100000;
            14'h0baa: o_data_a = 16'b1110001100001000;
            14'h0bab: o_data_a = 16'b0000000000000011;
            14'h0bac: o_data_a = 16'b1111110111100000;
            14'h0bad: o_data_a = 16'b1110110111100000;
            14'h0bae: o_data_a = 16'b1111110000010000;
            14'h0baf: o_data_a = 16'b0000000000000000;
            14'h0bb0: o_data_a = 16'b1111110111101000;
            14'h0bb1: o_data_a = 16'b1110110010100000;
            14'h0bb2: o_data_a = 16'b1110001100001000;
            14'h0bb3: o_data_a = 16'b0000000000000000;
            14'h0bb4: o_data_a = 16'b1111110010101000;
            14'h0bb5: o_data_a = 16'b1111110000010000;
            14'h0bb6: o_data_a = 16'b1110110010100000;
            14'h0bb7: o_data_a = 16'b1111000010001000;
            14'h0bb8: o_data_a = 16'b0000000000000011;
            14'h0bb9: o_data_a = 16'b1111110111100000;
            14'h0bba: o_data_a = 16'b1111110000010000;
            14'h0bbb: o_data_a = 16'b0000000000000000;
            14'h0bbc: o_data_a = 16'b1111110111101000;
            14'h0bbd: o_data_a = 16'b1110110010100000;
            14'h0bbe: o_data_a = 16'b1110001100001000;
            14'h0bbf: o_data_a = 16'b0000000000000011;
            14'h0bc0: o_data_a = 16'b1111110000010000;
            14'h0bc1: o_data_a = 16'b0000000000000011;
            14'h0bc2: o_data_a = 16'b1110000010100000;
            14'h0bc3: o_data_a = 16'b1111110000010000;
            14'h0bc4: o_data_a = 16'b0000000000000000;
            14'h0bc5: o_data_a = 16'b1111110111101000;
            14'h0bc6: o_data_a = 16'b1110110010100000;
            14'h0bc7: o_data_a = 16'b1110001100001000;
            14'h0bc8: o_data_a = 16'b0000000000000000;
            14'h0bc9: o_data_a = 16'b1111110010101000;
            14'h0bca: o_data_a = 16'b1111110000010000;
            14'h0bcb: o_data_a = 16'b1110110010100000;
            14'h0bcc: o_data_a = 16'b1111000010001000;
            14'h0bcd: o_data_a = 16'b0000000000000100;
            14'h0bce: o_data_a = 16'b1110110000010000;
            14'h0bcf: o_data_a = 16'b0000000000001101;
            14'h0bd0: o_data_a = 16'b1110001100001000;
            14'h0bd1: o_data_a = 16'b0101011101010010;
            14'h0bd2: o_data_a = 16'b1110110000010000;
            14'h0bd3: o_data_a = 16'b0000000000001110;
            14'h0bd4: o_data_a = 16'b1110001100001000;
            14'h0bd5: o_data_a = 16'b0000101111011001;
            14'h0bd6: o_data_a = 16'b1110110000010000;
            14'h0bd7: o_data_a = 16'b0000000001011111;
            14'h0bd8: o_data_a = 16'b1110101010000111;
            14'h0bd9: o_data_a = 16'b0000000000000000;
            14'h0bda: o_data_a = 16'b1111110010101000;
            14'h0bdb: o_data_a = 16'b1111110000010000;
            14'h0bdc: o_data_a = 16'b0000000000000101;
            14'h0bdd: o_data_a = 16'b1110001100001000;
            14'h0bde: o_data_a = 16'b0000000000000000;
            14'h0bdf: o_data_a = 16'b1111110111001000;
            14'h0be0: o_data_a = 16'b1111110010100000;
            14'h0be1: o_data_a = 16'b1110101010001000;
            14'h0be2: o_data_a = 16'b0000000000110110;
            14'h0be3: o_data_a = 16'b1110101010000111;
            14'h0be4: o_data_a = 16'b0000000000000010;
            14'h0be5: o_data_a = 16'b1111110000100000;
            14'h0be6: o_data_a = 16'b1111110000010000;
            14'h0be7: o_data_a = 16'b0000000000000000;
            14'h0be8: o_data_a = 16'b1111110111101000;
            14'h0be9: o_data_a = 16'b1110110010100000;
            14'h0bea: o_data_a = 16'b1110001100001000;
            14'h0beb: o_data_a = 16'b0000000000000000;
            14'h0bec: o_data_a = 16'b1111110010101000;
            14'h0bed: o_data_a = 16'b1111110000010000;
            14'h0bee: o_data_a = 16'b0000000000000011;
            14'h0bef: o_data_a = 16'b1110001100001000;
            14'h0bf0: o_data_a = 16'b0000000000000010;
            14'h0bf1: o_data_a = 16'b1111110111100000;
            14'h0bf2: o_data_a = 16'b1111110000010000;
            14'h0bf3: o_data_a = 16'b0000000000000000;
            14'h0bf4: o_data_a = 16'b1111110111101000;
            14'h0bf5: o_data_a = 16'b1110110010100000;
            14'h0bf6: o_data_a = 16'b1110001100001000;
            14'h0bf7: o_data_a = 16'b0000000000000000;
            14'h0bf8: o_data_a = 16'b1111110010101000;
            14'h0bf9: o_data_a = 16'b1111110000010000;
            14'h0bfa: o_data_a = 16'b0000000000000011;
            14'h0bfb: o_data_a = 16'b1111110111100000;
            14'h0bfc: o_data_a = 16'b1110110111100000;
            14'h0bfd: o_data_a = 16'b1110110111100000;
            14'h0bfe: o_data_a = 16'b1110110111100000;
            14'h0bff: o_data_a = 16'b1110001100001000;
            14'h0c00: o_data_a = 16'b0000000000000000;
            14'h0c01: o_data_a = 16'b1111110111001000;
            14'h0c02: o_data_a = 16'b1111110010100000;
            14'h0c03: o_data_a = 16'b1110101010001000;
            14'h0c04: o_data_a = 16'b0000000000110110;
            14'h0c05: o_data_a = 16'b1110101010000111;
            14'h0c06: o_data_a = 16'b0000000000000010;
            14'h0c07: o_data_a = 16'b1111110000100000;
            14'h0c08: o_data_a = 16'b1111110000010000;
            14'h0c09: o_data_a = 16'b0000000000000000;
            14'h0c0a: o_data_a = 16'b1111110111101000;
            14'h0c0b: o_data_a = 16'b1110110010100000;
            14'h0c0c: o_data_a = 16'b1110001100001000;
            14'h0c0d: o_data_a = 16'b0000000000000000;
            14'h0c0e: o_data_a = 16'b1111110010101000;
            14'h0c0f: o_data_a = 16'b1111110000010000;
            14'h0c10: o_data_a = 16'b0000000000000011;
            14'h0c11: o_data_a = 16'b1110001100001000;
            14'h0c12: o_data_a = 16'b0000000000000011;
            14'h0c13: o_data_a = 16'b1111110000100000;
            14'h0c14: o_data_a = 16'b1111110000010000;
            14'h0c15: o_data_a = 16'b0000000000000000;
            14'h0c16: o_data_a = 16'b1111110111101000;
            14'h0c17: o_data_a = 16'b1110110010100000;
            14'h0c18: o_data_a = 16'b1110001100001000;
            14'h0c19: o_data_a = 16'b0000000000110110;
            14'h0c1a: o_data_a = 16'b1110101010000111;
            14'h0c1b: o_data_a = 16'b0000000000000010;
            14'h0c1c: o_data_a = 16'b1111110000100000;
            14'h0c1d: o_data_a = 16'b1111110000010000;
            14'h0c1e: o_data_a = 16'b0000000000000000;
            14'h0c1f: o_data_a = 16'b1111110111101000;
            14'h0c20: o_data_a = 16'b1110110010100000;
            14'h0c21: o_data_a = 16'b1110001100001000;
            14'h0c22: o_data_a = 16'b0000000000000000;
            14'h0c23: o_data_a = 16'b1111110010101000;
            14'h0c24: o_data_a = 16'b1111110000010000;
            14'h0c25: o_data_a = 16'b0000000000000011;
            14'h0c26: o_data_a = 16'b1110001100001000;
            14'h0c27: o_data_a = 16'b0000000000000011;
            14'h0c28: o_data_a = 16'b1111110000100000;
            14'h0c29: o_data_a = 16'b1111110000010000;
            14'h0c2a: o_data_a = 16'b0000000000000000;
            14'h0c2b: o_data_a = 16'b1111110111101000;
            14'h0c2c: o_data_a = 16'b1110110010100000;
            14'h0c2d: o_data_a = 16'b1110001100001000;
            14'h0c2e: o_data_a = 16'b0000000000000011;
            14'h0c2f: o_data_a = 16'b1111110111100000;
            14'h0c30: o_data_a = 16'b1110110111100000;
            14'h0c31: o_data_a = 16'b1111110000010000;
            14'h0c32: o_data_a = 16'b0000000000000000;
            14'h0c33: o_data_a = 16'b1111110111101000;
            14'h0c34: o_data_a = 16'b1110110010100000;
            14'h0c35: o_data_a = 16'b1110001100001000;
            14'h0c36: o_data_a = 16'b0000000000000000;
            14'h0c37: o_data_a = 16'b1111110010101000;
            14'h0c38: o_data_a = 16'b1111110000010000;
            14'h0c39: o_data_a = 16'b1110110010100000;
            14'h0c3a: o_data_a = 16'b1111000010001000;
            14'h0c3b: o_data_a = 16'b0000000000110110;
            14'h0c3c: o_data_a = 16'b1110101010000111;
            14'h0c3d: o_data_a = 16'b0000000000000010;
            14'h0c3e: o_data_a = 16'b1111110000100000;
            14'h0c3f: o_data_a = 16'b1111110000010000;
            14'h0c40: o_data_a = 16'b0000000000000000;
            14'h0c41: o_data_a = 16'b1111110111101000;
            14'h0c42: o_data_a = 16'b1110110010100000;
            14'h0c43: o_data_a = 16'b1110001100001000;
            14'h0c44: o_data_a = 16'b0000000000000000;
            14'h0c45: o_data_a = 16'b1111110010101000;
            14'h0c46: o_data_a = 16'b1111110000010000;
            14'h0c47: o_data_a = 16'b0000000000000011;
            14'h0c48: o_data_a = 16'b1110001100001000;
            14'h0c49: o_data_a = 16'b0000000000000011;
            14'h0c4a: o_data_a = 16'b1111110000010000;
            14'h0c4b: o_data_a = 16'b0000000000000000;
            14'h0c4c: o_data_a = 16'b1111110111101000;
            14'h0c4d: o_data_a = 16'b1110110010100000;
            14'h0c4e: o_data_a = 16'b1110001100001000;
            14'h0c4f: o_data_a = 16'b0000000000000001;
            14'h0c50: o_data_a = 16'b1110110000010000;
            14'h0c51: o_data_a = 16'b0000000000001101;
            14'h0c52: o_data_a = 16'b1110001100001000;
            14'h0c53: o_data_a = 16'b0000101101001100;
            14'h0c54: o_data_a = 16'b1110110000010000;
            14'h0c55: o_data_a = 16'b0000000000001110;
            14'h0c56: o_data_a = 16'b1110001100001000;
            14'h0c57: o_data_a = 16'b0000110001011011;
            14'h0c58: o_data_a = 16'b1110110000010000;
            14'h0c59: o_data_a = 16'b0000000001011111;
            14'h0c5a: o_data_a = 16'b1110101010000111;
            14'h0c5b: o_data_a = 16'b0000000000000000;
            14'h0c5c: o_data_a = 16'b1111110010101000;
            14'h0c5d: o_data_a = 16'b1111110000010000;
            14'h0c5e: o_data_a = 16'b0000000000000101;
            14'h0c5f: o_data_a = 16'b1110001100001000;
            14'h0c60: o_data_a = 16'b0000000000000010;
            14'h0c61: o_data_a = 16'b1111110111100000;
            14'h0c62: o_data_a = 16'b1111110000010000;
            14'h0c63: o_data_a = 16'b0000000000000000;
            14'h0c64: o_data_a = 16'b1111110111101000;
            14'h0c65: o_data_a = 16'b1110110010100000;
            14'h0c66: o_data_a = 16'b1110001100001000;
            14'h0c67: o_data_a = 16'b0000000000000000;
            14'h0c68: o_data_a = 16'b1111110010101000;
            14'h0c69: o_data_a = 16'b1111110000010000;
            14'h0c6a: o_data_a = 16'b0000000000000011;
            14'h0c6b: o_data_a = 16'b1111110111100000;
            14'h0c6c: o_data_a = 16'b1110110111100000;
            14'h0c6d: o_data_a = 16'b1110001100001000;
            14'h0c6e: o_data_a = 16'b0000000000000011;
            14'h0c6f: o_data_a = 16'b1111110000010000;
            14'h0c70: o_data_a = 16'b0000000000000000;
            14'h0c71: o_data_a = 16'b1111110111101000;
            14'h0c72: o_data_a = 16'b1110110010100000;
            14'h0c73: o_data_a = 16'b1110001100001000;
            14'h0c74: o_data_a = 16'b0000000000000001;
            14'h0c75: o_data_a = 16'b1110110000010000;
            14'h0c76: o_data_a = 16'b0000000000001101;
            14'h0c77: o_data_a = 16'b1110001100001000;
            14'h0c78: o_data_a = 16'b0000101100001011;
            14'h0c79: o_data_a = 16'b1110110000010000;
            14'h0c7a: o_data_a = 16'b0000000000001110;
            14'h0c7b: o_data_a = 16'b1110001100001000;
            14'h0c7c: o_data_a = 16'b0000110010000000;
            14'h0c7d: o_data_a = 16'b1110110000010000;
            14'h0c7e: o_data_a = 16'b0000000001011111;
            14'h0c7f: o_data_a = 16'b1110101010000111;
            14'h0c80: o_data_a = 16'b0000000000000000;
            14'h0c81: o_data_a = 16'b1111110010101000;
            14'h0c82: o_data_a = 16'b1111110000010000;
            14'h0c83: o_data_a = 16'b0000000000000101;
            14'h0c84: o_data_a = 16'b1110001100001000;
            14'h0c85: o_data_a = 16'b0000000000000000;
            14'h0c86: o_data_a = 16'b1111110111001000;
            14'h0c87: o_data_a = 16'b1111110010100000;
            14'h0c88: o_data_a = 16'b1110101010001000;
            14'h0c89: o_data_a = 16'b0000000000110110;
            14'h0c8a: o_data_a = 16'b1110101010000111;
            14'h0c8b: o_data_a = 16'b0000000000000010;
            14'h0c8c: o_data_a = 16'b1111110000100000;
            14'h0c8d: o_data_a = 16'b1111110000010000;
            14'h0c8e: o_data_a = 16'b0000000000000000;
            14'h0c8f: o_data_a = 16'b1111110111101000;
            14'h0c90: o_data_a = 16'b1110110010100000;
            14'h0c91: o_data_a = 16'b1110001100001000;
            14'h0c92: o_data_a = 16'b0000000000000000;
            14'h0c93: o_data_a = 16'b1111110010101000;
            14'h0c94: o_data_a = 16'b1111110000010000;
            14'h0c95: o_data_a = 16'b0000000000000011;
            14'h0c96: o_data_a = 16'b1110001100001000;
            14'h0c97: o_data_a = 16'b0000000000000011;
            14'h0c98: o_data_a = 16'b1111110000010000;
            14'h0c99: o_data_a = 16'b0000000000000100;
            14'h0c9a: o_data_a = 16'b1110000010100000;
            14'h0c9b: o_data_a = 16'b1111110000010000;
            14'h0c9c: o_data_a = 16'b0000000000000000;
            14'h0c9d: o_data_a = 16'b1111110111101000;
            14'h0c9e: o_data_a = 16'b1110110010100000;
            14'h0c9f: o_data_a = 16'b1110001100001000;
            14'h0ca0: o_data_a = 16'b0000000000000000;
            14'h0ca1: o_data_a = 16'b1111110111001000;
            14'h0ca2: o_data_a = 16'b1111110010100000;
            14'h0ca3: o_data_a = 16'b1110111111001000;
            14'h0ca4: o_data_a = 16'b0000110010101000;
            14'h0ca5: o_data_a = 16'b1110110000010000;
            14'h0ca6: o_data_a = 16'b0000000000000110;
            14'h0ca7: o_data_a = 16'b1110101010000111;
            14'h0ca8: o_data_a = 16'b0000000000000000;
            14'h0ca9: o_data_a = 16'b1111110010101000;
            14'h0caa: o_data_a = 16'b1111110000010000;
            14'h0cab: o_data_a = 16'b0000110010101111;
            14'h0cac: o_data_a = 16'b1110001100000101;
            14'h0cad: o_data_a = 16'b0000110111000101;
            14'h0cae: o_data_a = 16'b1110101010000111;
            14'h0caf: o_data_a = 16'b0000000000000011;
            14'h0cb0: o_data_a = 16'b1111110000100000;
            14'h0cb1: o_data_a = 16'b1111110000010000;
            14'h0cb2: o_data_a = 16'b0000000000000000;
            14'h0cb3: o_data_a = 16'b1111110111101000;
            14'h0cb4: o_data_a = 16'b1110110010100000;
            14'h0cb5: o_data_a = 16'b1110001100001000;
            14'h0cb6: o_data_a = 16'b0000000000000100;
            14'h0cb7: o_data_a = 16'b1110110000010000;
            14'h0cb8: o_data_a = 16'b0000000000000000;
            14'h0cb9: o_data_a = 16'b1111110111101000;
            14'h0cba: o_data_a = 16'b1110110010100000;
            14'h0cbb: o_data_a = 16'b1110001100001000;
            14'h0cbc: o_data_a = 16'b0000000000000000;
            14'h0cbd: o_data_a = 16'b1111110010101000;
            14'h0cbe: o_data_a = 16'b1111110000010000;
            14'h0cbf: o_data_a = 16'b1110110010100000;
            14'h0cc0: o_data_a = 16'b1111000111001000;
            14'h0cc1: o_data_a = 16'b0000000000000000;
            14'h0cc2: o_data_a = 16'b1111110010101000;
            14'h0cc3: o_data_a = 16'b1111110000010000;
            14'h0cc4: o_data_a = 16'b0000000000000011;
            14'h0cc5: o_data_a = 16'b1111110000100000;
            14'h0cc6: o_data_a = 16'b1110001100001000;
            14'h0cc7: o_data_a = 16'b0000000000000011;
            14'h0cc8: o_data_a = 16'b1111110000100000;
            14'h0cc9: o_data_a = 16'b1111110000010000;
            14'h0cca: o_data_a = 16'b0000000000000000;
            14'h0ccb: o_data_a = 16'b1111110111101000;
            14'h0ccc: o_data_a = 16'b1110110010100000;
            14'h0ccd: o_data_a = 16'b1110001100001000;
            14'h0cce: o_data_a = 16'b0000000000000000;
            14'h0ccf: o_data_a = 16'b1111110111001000;
            14'h0cd0: o_data_a = 16'b1111110010100000;
            14'h0cd1: o_data_a = 16'b1110101010001000;
            14'h0cd2: o_data_a = 16'b0000110011010110;
            14'h0cd3: o_data_a = 16'b1110110000010000;
            14'h0cd4: o_data_a = 16'b0000000000100110;
            14'h0cd5: o_data_a = 16'b1110101010000111;
            14'h0cd6: o_data_a = 16'b0000000000000000;
            14'h0cd7: o_data_a = 16'b1111110010101000;
            14'h0cd8: o_data_a = 16'b1111110000010000;
            14'h0cd9: o_data_a = 16'b0000110011011101;
            14'h0cda: o_data_a = 16'b1110001100000101;
            14'h0cdb: o_data_a = 16'b0000110011100111;
            14'h0cdc: o_data_a = 16'b1110101010000111;
            14'h0cdd: o_data_a = 16'b0000000000000000;
            14'h0cde: o_data_a = 16'b1111110111001000;
            14'h0cdf: o_data_a = 16'b1111110010100000;
            14'h0ce0: o_data_a = 16'b1110101010001000;
            14'h0ce1: o_data_a = 16'b0000000000000000;
            14'h0ce2: o_data_a = 16'b1111110010101000;
            14'h0ce3: o_data_a = 16'b1111110000010000;
            14'h0ce4: o_data_a = 16'b0000000000000011;
            14'h0ce5: o_data_a = 16'b1111110000100000;
            14'h0ce6: o_data_a = 16'b1110001100001000;
            14'h0ce7: o_data_a = 16'b0000000000000000;
            14'h0ce8: o_data_a = 16'b1111110111001000;
            14'h0ce9: o_data_a = 16'b1111110010100000;
            14'h0cea: o_data_a = 16'b1110101010001000;
            14'h0ceb: o_data_a = 16'b0000000000000001;
            14'h0cec: o_data_a = 16'b1110110000010000;
            14'h0ced: o_data_a = 16'b0000000000001101;
            14'h0cee: o_data_a = 16'b1110001100001000;
            14'h0cef: o_data_a = 16'b0101000110011001;
            14'h0cf0: o_data_a = 16'b1110110000010000;
            14'h0cf1: o_data_a = 16'b0000000000001110;
            14'h0cf2: o_data_a = 16'b1110001100001000;
            14'h0cf3: o_data_a = 16'b0000110011110111;
            14'h0cf4: o_data_a = 16'b1110110000010000;
            14'h0cf5: o_data_a = 16'b0000000001011111;
            14'h0cf6: o_data_a = 16'b1110101010000111;
            14'h0cf7: o_data_a = 16'b0000000000000000;
            14'h0cf8: o_data_a = 16'b1111110010101000;
            14'h0cf9: o_data_a = 16'b1111110000010000;
            14'h0cfa: o_data_a = 16'b0000000000000101;
            14'h0cfb: o_data_a = 16'b1110001100001000;
            14'h0cfc: o_data_a = 16'b0000000000000011;
            14'h0cfd: o_data_a = 16'b1111110000100000;
            14'h0cfe: o_data_a = 16'b1111110000010000;
            14'h0cff: o_data_a = 16'b0000000000000000;
            14'h0d00: o_data_a = 16'b1111110111101000;
            14'h0d01: o_data_a = 16'b1110110010100000;
            14'h0d02: o_data_a = 16'b1110001100001000;
            14'h0d03: o_data_a = 16'b0000000000000011;
            14'h0d04: o_data_a = 16'b1111110111100000;
            14'h0d05: o_data_a = 16'b1110110111100000;
            14'h0d06: o_data_a = 16'b1111110000010000;
            14'h0d07: o_data_a = 16'b0000000000000000;
            14'h0d08: o_data_a = 16'b1111110111101000;
            14'h0d09: o_data_a = 16'b1110110010100000;
            14'h0d0a: o_data_a = 16'b1110001100001000;
            14'h0d0b: o_data_a = 16'b0000000000000000;
            14'h0d0c: o_data_a = 16'b1111110010101000;
            14'h0d0d: o_data_a = 16'b1111110000010000;
            14'h0d0e: o_data_a = 16'b1110110010100000;
            14'h0d0f: o_data_a = 16'b1111000010001000;
            14'h0d10: o_data_a = 16'b0000000000000000;
            14'h0d11: o_data_a = 16'b1111110111001000;
            14'h0d12: o_data_a = 16'b1111110010100000;
            14'h0d13: o_data_a = 16'b1110111111001000;
            14'h0d14: o_data_a = 16'b0000000000000000;
            14'h0d15: o_data_a = 16'b1111110010101000;
            14'h0d16: o_data_a = 16'b1111110000010000;
            14'h0d17: o_data_a = 16'b1110110010100000;
            14'h0d18: o_data_a = 16'b1111000010001000;
            14'h0d19: o_data_a = 16'b0000000000000011;
            14'h0d1a: o_data_a = 16'b1111110111100000;
            14'h0d1b: o_data_a = 16'b1111110000010000;
            14'h0d1c: o_data_a = 16'b0000000000000000;
            14'h0d1d: o_data_a = 16'b1111110111101000;
            14'h0d1e: o_data_a = 16'b1110110010100000;
            14'h0d1f: o_data_a = 16'b1110001100001000;
            14'h0d20: o_data_a = 16'b0000000000000011;
            14'h0d21: o_data_a = 16'b1111110000100000;
            14'h0d22: o_data_a = 16'b1111110000010000;
            14'h0d23: o_data_a = 16'b0000000000000000;
            14'h0d24: o_data_a = 16'b1111110111101000;
            14'h0d25: o_data_a = 16'b1110110010100000;
            14'h0d26: o_data_a = 16'b1110001100001000;
            14'h0d27: o_data_a = 16'b0000000000000011;
            14'h0d28: o_data_a = 16'b1111110111100000;
            14'h0d29: o_data_a = 16'b1110110111100000;
            14'h0d2a: o_data_a = 16'b1111110000010000;
            14'h0d2b: o_data_a = 16'b0000000000000000;
            14'h0d2c: o_data_a = 16'b1111110111101000;
            14'h0d2d: o_data_a = 16'b1110110010100000;
            14'h0d2e: o_data_a = 16'b1110001100001000;
            14'h0d2f: o_data_a = 16'b0000000000000000;
            14'h0d30: o_data_a = 16'b1111110010101000;
            14'h0d31: o_data_a = 16'b1111110000010000;
            14'h0d32: o_data_a = 16'b1110110010100000;
            14'h0d33: o_data_a = 16'b1111000010001000;
            14'h0d34: o_data_a = 16'b0000000000000100;
            14'h0d35: o_data_a = 16'b1110110000010000;
            14'h0d36: o_data_a = 16'b0000000000000000;
            14'h0d37: o_data_a = 16'b1111110111101000;
            14'h0d38: o_data_a = 16'b1110110010100000;
            14'h0d39: o_data_a = 16'b1110001100001000;
            14'h0d3a: o_data_a = 16'b0000000000000000;
            14'h0d3b: o_data_a = 16'b1111110010101000;
            14'h0d3c: o_data_a = 16'b1111110000010000;
            14'h0d3d: o_data_a = 16'b1110110010100000;
            14'h0d3e: o_data_a = 16'b1111000010001000;
            14'h0d3f: o_data_a = 16'b0000000000000011;
            14'h0d40: o_data_a = 16'b1111110111100000;
            14'h0d41: o_data_a = 16'b1111110000010000;
            14'h0d42: o_data_a = 16'b0000000000000000;
            14'h0d43: o_data_a = 16'b1111110111101000;
            14'h0d44: o_data_a = 16'b1110110010100000;
            14'h0d45: o_data_a = 16'b1110001100001000;
            14'h0d46: o_data_a = 16'b0000000000000011;
            14'h0d47: o_data_a = 16'b1111110000010000;
            14'h0d48: o_data_a = 16'b0000000000000011;
            14'h0d49: o_data_a = 16'b1110000010100000;
            14'h0d4a: o_data_a = 16'b1111110000010000;
            14'h0d4b: o_data_a = 16'b0000000000000000;
            14'h0d4c: o_data_a = 16'b1111110111101000;
            14'h0d4d: o_data_a = 16'b1110110010100000;
            14'h0d4e: o_data_a = 16'b1110001100001000;
            14'h0d4f: o_data_a = 16'b0000000000000000;
            14'h0d50: o_data_a = 16'b1111110010101000;
            14'h0d51: o_data_a = 16'b1111110000010000;
            14'h0d52: o_data_a = 16'b1110110010100000;
            14'h0d53: o_data_a = 16'b1111000010001000;
            14'h0d54: o_data_a = 16'b0000000000000100;
            14'h0d55: o_data_a = 16'b1110110000010000;
            14'h0d56: o_data_a = 16'b0000000000001101;
            14'h0d57: o_data_a = 16'b1110001100001000;
            14'h0d58: o_data_a = 16'b0101011101010010;
            14'h0d59: o_data_a = 16'b1110110000010000;
            14'h0d5a: o_data_a = 16'b0000000000001110;
            14'h0d5b: o_data_a = 16'b1110001100001000;
            14'h0d5c: o_data_a = 16'b0000110101100000;
            14'h0d5d: o_data_a = 16'b1110110000010000;
            14'h0d5e: o_data_a = 16'b0000000001011111;
            14'h0d5f: o_data_a = 16'b1110101010000111;
            14'h0d60: o_data_a = 16'b0000000000000000;
            14'h0d61: o_data_a = 16'b1111110010101000;
            14'h0d62: o_data_a = 16'b1111110000010000;
            14'h0d63: o_data_a = 16'b0000000000000101;
            14'h0d64: o_data_a = 16'b1110001100001000;
            14'h0d65: o_data_a = 16'b0000000000000000;
            14'h0d66: o_data_a = 16'b1111110111001000;
            14'h0d67: o_data_a = 16'b1111110010100000;
            14'h0d68: o_data_a = 16'b1110101010001000;
            14'h0d69: o_data_a = 16'b0000000000000000;
            14'h0d6a: o_data_a = 16'b1111110010100000;
            14'h0d6b: o_data_a = 16'b1111110001001000;
            14'h0d6c: o_data_a = 16'b0000000000000001;
            14'h0d6d: o_data_a = 16'b1110110000010000;
            14'h0d6e: o_data_a = 16'b0000000000001101;
            14'h0d6f: o_data_a = 16'b1110001100001000;
            14'h0d70: o_data_a = 16'b0101000110011001;
            14'h0d71: o_data_a = 16'b1110110000010000;
            14'h0d72: o_data_a = 16'b0000000000001110;
            14'h0d73: o_data_a = 16'b1110001100001000;
            14'h0d74: o_data_a = 16'b0000110101111000;
            14'h0d75: o_data_a = 16'b1110110000010000;
            14'h0d76: o_data_a = 16'b0000000001011111;
            14'h0d77: o_data_a = 16'b1110101010000111;
            14'h0d78: o_data_a = 16'b0000000000000000;
            14'h0d79: o_data_a = 16'b1111110010101000;
            14'h0d7a: o_data_a = 16'b1111110000010000;
            14'h0d7b: o_data_a = 16'b0000000000000101;
            14'h0d7c: o_data_a = 16'b1110001100001000;
            14'h0d7d: o_data_a = 16'b0000000000000011;
            14'h0d7e: o_data_a = 16'b1111110000100000;
            14'h0d7f: o_data_a = 16'b1111110000010000;
            14'h0d80: o_data_a = 16'b0000000000000000;
            14'h0d81: o_data_a = 16'b1111110111101000;
            14'h0d82: o_data_a = 16'b1110110010100000;
            14'h0d83: o_data_a = 16'b1110001100001000;
            14'h0d84: o_data_a = 16'b0000000000000011;
            14'h0d85: o_data_a = 16'b1111110111100000;
            14'h0d86: o_data_a = 16'b1111110000010000;
            14'h0d87: o_data_a = 16'b0000000000000000;
            14'h0d88: o_data_a = 16'b1111110111101000;
            14'h0d89: o_data_a = 16'b1110110010100000;
            14'h0d8a: o_data_a = 16'b1110001100001000;
            14'h0d8b: o_data_a = 16'b0000000000000011;
            14'h0d8c: o_data_a = 16'b1111110000100000;
            14'h0d8d: o_data_a = 16'b1111110000010000;
            14'h0d8e: o_data_a = 16'b0000000000000000;
            14'h0d8f: o_data_a = 16'b1111110111101000;
            14'h0d90: o_data_a = 16'b1110110010100000;
            14'h0d91: o_data_a = 16'b1110001100001000;
            14'h0d92: o_data_a = 16'b0000000000000011;
            14'h0d93: o_data_a = 16'b1110110000010000;
            14'h0d94: o_data_a = 16'b0000000000000000;
            14'h0d95: o_data_a = 16'b1111110111101000;
            14'h0d96: o_data_a = 16'b1110110010100000;
            14'h0d97: o_data_a = 16'b1110001100001000;
            14'h0d98: o_data_a = 16'b0000000000000000;
            14'h0d99: o_data_a = 16'b1111110010101000;
            14'h0d9a: o_data_a = 16'b1111110000010000;
            14'h0d9b: o_data_a = 16'b1110110010100000;
            14'h0d9c: o_data_a = 16'b1111000010001000;
            14'h0d9d: o_data_a = 16'b0000000000000011;
            14'h0d9e: o_data_a = 16'b1111110111100000;
            14'h0d9f: o_data_a = 16'b1111110000010000;
            14'h0da0: o_data_a = 16'b0000000000000000;
            14'h0da1: o_data_a = 16'b1111110111101000;
            14'h0da2: o_data_a = 16'b1110110010100000;
            14'h0da3: o_data_a = 16'b1110001100001000;
            14'h0da4: o_data_a = 16'b0000000000000011;
            14'h0da5: o_data_a = 16'b1111110000010000;
            14'h0da6: o_data_a = 16'b0000000000000011;
            14'h0da7: o_data_a = 16'b1110000010100000;
            14'h0da8: o_data_a = 16'b1111110000010000;
            14'h0da9: o_data_a = 16'b0000000000000000;
            14'h0daa: o_data_a = 16'b1111110111101000;
            14'h0dab: o_data_a = 16'b1110110010100000;
            14'h0dac: o_data_a = 16'b1110001100001000;
            14'h0dad: o_data_a = 16'b0000000000000000;
            14'h0dae: o_data_a = 16'b1111110010101000;
            14'h0daf: o_data_a = 16'b1111110000010000;
            14'h0db0: o_data_a = 16'b1110110010100000;
            14'h0db1: o_data_a = 16'b1111000010001000;
            14'h0db2: o_data_a = 16'b0000000000000100;
            14'h0db3: o_data_a = 16'b1110110000010000;
            14'h0db4: o_data_a = 16'b0000000000001101;
            14'h0db5: o_data_a = 16'b1110001100001000;
            14'h0db6: o_data_a = 16'b0101011101010010;
            14'h0db7: o_data_a = 16'b1110110000010000;
            14'h0db8: o_data_a = 16'b0000000000001110;
            14'h0db9: o_data_a = 16'b1110001100001000;
            14'h0dba: o_data_a = 16'b0000110110111110;
            14'h0dbb: o_data_a = 16'b1110110000010000;
            14'h0dbc: o_data_a = 16'b0000000001011111;
            14'h0dbd: o_data_a = 16'b1110101010000111;
            14'h0dbe: o_data_a = 16'b0000000000000000;
            14'h0dbf: o_data_a = 16'b1111110010101000;
            14'h0dc0: o_data_a = 16'b1111110000010000;
            14'h0dc1: o_data_a = 16'b0000000000000101;
            14'h0dc2: o_data_a = 16'b1110001100001000;
            14'h0dc3: o_data_a = 16'b0000111011110111;
            14'h0dc4: o_data_a = 16'b1110101010000111;
            14'h0dc5: o_data_a = 16'b0000000000000011;
            14'h0dc6: o_data_a = 16'b1111110000100000;
            14'h0dc7: o_data_a = 16'b1111110000010000;
            14'h0dc8: o_data_a = 16'b0000000000000000;
            14'h0dc9: o_data_a = 16'b1111110111101000;
            14'h0dca: o_data_a = 16'b1110110010100000;
            14'h0dcb: o_data_a = 16'b1110001100001000;
            14'h0dcc: o_data_a = 16'b0000000000000100;
            14'h0dcd: o_data_a = 16'b1110110000010000;
            14'h0dce: o_data_a = 16'b0000000000000000;
            14'h0dcf: o_data_a = 16'b1111110111101000;
            14'h0dd0: o_data_a = 16'b1110110010100000;
            14'h0dd1: o_data_a = 16'b1110001100001000;
            14'h0dd2: o_data_a = 16'b0000000000000000;
            14'h0dd3: o_data_a = 16'b1111110010101000;
            14'h0dd4: o_data_a = 16'b1111110000010000;
            14'h0dd5: o_data_a = 16'b1110110010100000;
            14'h0dd6: o_data_a = 16'b1111000010001000;
            14'h0dd7: o_data_a = 16'b0000000000000000;
            14'h0dd8: o_data_a = 16'b1111110010101000;
            14'h0dd9: o_data_a = 16'b1111110000010000;
            14'h0dda: o_data_a = 16'b0000000000000011;
            14'h0ddb: o_data_a = 16'b1111110000100000;
            14'h0ddc: o_data_a = 16'b1110001100001000;
            14'h0ddd: o_data_a = 16'b0000000000000011;
            14'h0dde: o_data_a = 16'b1111110000100000;
            14'h0ddf: o_data_a = 16'b1111110000010000;
            14'h0de0: o_data_a = 16'b0000000000000000;
            14'h0de1: o_data_a = 16'b1111110111101000;
            14'h0de2: o_data_a = 16'b1110110010100000;
            14'h0de3: o_data_a = 16'b1110001100001000;
            14'h0de4: o_data_a = 16'b0000000000000011;
            14'h0de5: o_data_a = 16'b1111110111100000;
            14'h0de6: o_data_a = 16'b1110110111100000;
            14'h0de7: o_data_a = 16'b1111110000010000;
            14'h0de8: o_data_a = 16'b0000000000000000;
            14'h0de9: o_data_a = 16'b1111110111101000;
            14'h0dea: o_data_a = 16'b1110110010100000;
            14'h0deb: o_data_a = 16'b1110001100001000;
            14'h0dec: o_data_a = 16'b0000000000000000;
            14'h0ded: o_data_a = 16'b1111110010101000;
            14'h0dee: o_data_a = 16'b1111110000010000;
            14'h0def: o_data_a = 16'b1110110010100000;
            14'h0df0: o_data_a = 16'b1111000010001000;
            14'h0df1: o_data_a = 16'b0000000111111111;
            14'h0df2: o_data_a = 16'b1110110000010000;
            14'h0df3: o_data_a = 16'b0000000000000000;
            14'h0df4: o_data_a = 16'b1111110111101000;
            14'h0df5: o_data_a = 16'b1110110010100000;
            14'h0df6: o_data_a = 16'b1110001100001000;
            14'h0df7: o_data_a = 16'b0000110111111011;
            14'h0df8: o_data_a = 16'b1110110000010000;
            14'h0df9: o_data_a = 16'b0000000000010110;
            14'h0dfa: o_data_a = 16'b1110101010000111;
            14'h0dfb: o_data_a = 16'b0000000000000000;
            14'h0dfc: o_data_a = 16'b1111110010101000;
            14'h0dfd: o_data_a = 16'b1111110000010000;
            14'h0dfe: o_data_a = 16'b0000111000000010;
            14'h0dff: o_data_a = 16'b1110001100000101;
            14'h0e00: o_data_a = 16'b0000111000011011;
            14'h0e01: o_data_a = 16'b1110101010000111;
            14'h0e02: o_data_a = 16'b0000000111111111;
            14'h0e03: o_data_a = 16'b1110110000010000;
            14'h0e04: o_data_a = 16'b0000000000000000;
            14'h0e05: o_data_a = 16'b1111110111101000;
            14'h0e06: o_data_a = 16'b1110110010100000;
            14'h0e07: o_data_a = 16'b1110001100001000;
            14'h0e08: o_data_a = 16'b0000000000000011;
            14'h0e09: o_data_a = 16'b1111110111100000;
            14'h0e0a: o_data_a = 16'b1110110111100000;
            14'h0e0b: o_data_a = 16'b1111110000010000;
            14'h0e0c: o_data_a = 16'b0000000000000000;
            14'h0e0d: o_data_a = 16'b1111110111101000;
            14'h0e0e: o_data_a = 16'b1110110010100000;
            14'h0e0f: o_data_a = 16'b1110001100001000;
            14'h0e10: o_data_a = 16'b0000000000000000;
            14'h0e11: o_data_a = 16'b1111110010101000;
            14'h0e12: o_data_a = 16'b1111110000010000;
            14'h0e13: o_data_a = 16'b1110110010100000;
            14'h0e14: o_data_a = 16'b1111000111001000;
            14'h0e15: o_data_a = 16'b0000000000000000;
            14'h0e16: o_data_a = 16'b1111110010101000;
            14'h0e17: o_data_a = 16'b1111110000010000;
            14'h0e18: o_data_a = 16'b0000000000000011;
            14'h0e19: o_data_a = 16'b1111110000100000;
            14'h0e1a: o_data_a = 16'b1110001100001000;
            14'h0e1b: o_data_a = 16'b0000000000000000;
            14'h0e1c: o_data_a = 16'b1111110111001000;
            14'h0e1d: o_data_a = 16'b1111110010100000;
            14'h0e1e: o_data_a = 16'b1110101010001000;
            14'h0e1f: o_data_a = 16'b0000000000000001;
            14'h0e20: o_data_a = 16'b1110110000010000;
            14'h0e21: o_data_a = 16'b0000000000001101;
            14'h0e22: o_data_a = 16'b1110001100001000;
            14'h0e23: o_data_a = 16'b0101000110011001;
            14'h0e24: o_data_a = 16'b1110110000010000;
            14'h0e25: o_data_a = 16'b0000000000001110;
            14'h0e26: o_data_a = 16'b1110001100001000;
            14'h0e27: o_data_a = 16'b0000111000101011;
            14'h0e28: o_data_a = 16'b1110110000010000;
            14'h0e29: o_data_a = 16'b0000000001011111;
            14'h0e2a: o_data_a = 16'b1110101010000111;
            14'h0e2b: o_data_a = 16'b0000000000000000;
            14'h0e2c: o_data_a = 16'b1111110010101000;
            14'h0e2d: o_data_a = 16'b1111110000010000;
            14'h0e2e: o_data_a = 16'b0000000000000101;
            14'h0e2f: o_data_a = 16'b1110001100001000;
            14'h0e30: o_data_a = 16'b0000000000000011;
            14'h0e31: o_data_a = 16'b1111110000100000;
            14'h0e32: o_data_a = 16'b1111110000010000;
            14'h0e33: o_data_a = 16'b0000000000000000;
            14'h0e34: o_data_a = 16'b1111110111101000;
            14'h0e35: o_data_a = 16'b1110110010100000;
            14'h0e36: o_data_a = 16'b1110001100001000;
            14'h0e37: o_data_a = 16'b0000000000000100;
            14'h0e38: o_data_a = 16'b1110110000010000;
            14'h0e39: o_data_a = 16'b0000000000000000;
            14'h0e3a: o_data_a = 16'b1111110111101000;
            14'h0e3b: o_data_a = 16'b1110110010100000;
            14'h0e3c: o_data_a = 16'b1110001100001000;
            14'h0e3d: o_data_a = 16'b0000000000000000;
            14'h0e3e: o_data_a = 16'b1111110010101000;
            14'h0e3f: o_data_a = 16'b1111110000010000;
            14'h0e40: o_data_a = 16'b1110110010100000;
            14'h0e41: o_data_a = 16'b1111000111001000;
            14'h0e42: o_data_a = 16'b0000000000000011;
            14'h0e43: o_data_a = 16'b1111110111100000;
            14'h0e44: o_data_a = 16'b1111110000010000;
            14'h0e45: o_data_a = 16'b0000000000000000;
            14'h0e46: o_data_a = 16'b1111110111101000;
            14'h0e47: o_data_a = 16'b1110110010100000;
            14'h0e48: o_data_a = 16'b1110001100001000;
            14'h0e49: o_data_a = 16'b0000000000000011;
            14'h0e4a: o_data_a = 16'b1111110000100000;
            14'h0e4b: o_data_a = 16'b1111110000010000;
            14'h0e4c: o_data_a = 16'b0000000000000000;
            14'h0e4d: o_data_a = 16'b1111110111101000;
            14'h0e4e: o_data_a = 16'b1110110010100000;
            14'h0e4f: o_data_a = 16'b1110001100001000;
            14'h0e50: o_data_a = 16'b0000000000000000;
            14'h0e51: o_data_a = 16'b1111110111001000;
            14'h0e52: o_data_a = 16'b1111110010100000;
            14'h0e53: o_data_a = 16'b1110111111001000;
            14'h0e54: o_data_a = 16'b0000000000000000;
            14'h0e55: o_data_a = 16'b1111110010101000;
            14'h0e56: o_data_a = 16'b1111110000010000;
            14'h0e57: o_data_a = 16'b1110110010100000;
            14'h0e58: o_data_a = 16'b1111000111001000;
            14'h0e59: o_data_a = 16'b0000000000000011;
            14'h0e5a: o_data_a = 16'b1111110111100000;
            14'h0e5b: o_data_a = 16'b1111110000010000;
            14'h0e5c: o_data_a = 16'b0000000000000000;
            14'h0e5d: o_data_a = 16'b1111110111101000;
            14'h0e5e: o_data_a = 16'b1110110010100000;
            14'h0e5f: o_data_a = 16'b1110001100001000;
            14'h0e60: o_data_a = 16'b0000000000000011;
            14'h0e61: o_data_a = 16'b1111110000010000;
            14'h0e62: o_data_a = 16'b0000000000000011;
            14'h0e63: o_data_a = 16'b1110000010100000;
            14'h0e64: o_data_a = 16'b1111110000010000;
            14'h0e65: o_data_a = 16'b0000000000000000;
            14'h0e66: o_data_a = 16'b1111110111101000;
            14'h0e67: o_data_a = 16'b1110110010100000;
            14'h0e68: o_data_a = 16'b1110001100001000;
            14'h0e69: o_data_a = 16'b0000000000000000;
            14'h0e6a: o_data_a = 16'b1111110010101000;
            14'h0e6b: o_data_a = 16'b1111110000010000;
            14'h0e6c: o_data_a = 16'b1110110010100000;
            14'h0e6d: o_data_a = 16'b1111000010001000;
            14'h0e6e: o_data_a = 16'b0000000000000100;
            14'h0e6f: o_data_a = 16'b1110110000010000;
            14'h0e70: o_data_a = 16'b0000000000001101;
            14'h0e71: o_data_a = 16'b1110001100001000;
            14'h0e72: o_data_a = 16'b0101011101010010;
            14'h0e73: o_data_a = 16'b1110110000010000;
            14'h0e74: o_data_a = 16'b0000000000001110;
            14'h0e75: o_data_a = 16'b1110001100001000;
            14'h0e76: o_data_a = 16'b0000111001111010;
            14'h0e77: o_data_a = 16'b1110110000010000;
            14'h0e78: o_data_a = 16'b0000000001011111;
            14'h0e79: o_data_a = 16'b1110101010000111;
            14'h0e7a: o_data_a = 16'b0000000000000000;
            14'h0e7b: o_data_a = 16'b1111110010101000;
            14'h0e7c: o_data_a = 16'b1111110000010000;
            14'h0e7d: o_data_a = 16'b0000000000000101;
            14'h0e7e: o_data_a = 16'b1110001100001000;
            14'h0e7f: o_data_a = 16'b0000000000000000;
            14'h0e80: o_data_a = 16'b1111110111001000;
            14'h0e81: o_data_a = 16'b1111110010100000;
            14'h0e82: o_data_a = 16'b1110101010001000;
            14'h0e83: o_data_a = 16'b0000000000000000;
            14'h0e84: o_data_a = 16'b1111110010100000;
            14'h0e85: o_data_a = 16'b1111110001001000;
            14'h0e86: o_data_a = 16'b0000000000000001;
            14'h0e87: o_data_a = 16'b1110110000010000;
            14'h0e88: o_data_a = 16'b0000000000001101;
            14'h0e89: o_data_a = 16'b1110001100001000;
            14'h0e8a: o_data_a = 16'b0101000110011001;
            14'h0e8b: o_data_a = 16'b1110110000010000;
            14'h0e8c: o_data_a = 16'b0000000000001110;
            14'h0e8d: o_data_a = 16'b1110001100001000;
            14'h0e8e: o_data_a = 16'b0000111010010010;
            14'h0e8f: o_data_a = 16'b1110110000010000;
            14'h0e90: o_data_a = 16'b0000000001011111;
            14'h0e91: o_data_a = 16'b1110101010000111;
            14'h0e92: o_data_a = 16'b0000000000000000;
            14'h0e93: o_data_a = 16'b1111110010101000;
            14'h0e94: o_data_a = 16'b1111110000010000;
            14'h0e95: o_data_a = 16'b0000000000000101;
            14'h0e96: o_data_a = 16'b1110001100001000;
            14'h0e97: o_data_a = 16'b0000000000000011;
            14'h0e98: o_data_a = 16'b1111110000100000;
            14'h0e99: o_data_a = 16'b1111110000010000;
            14'h0e9a: o_data_a = 16'b0000000000000000;
            14'h0e9b: o_data_a = 16'b1111110111101000;
            14'h0e9c: o_data_a = 16'b1110110010100000;
            14'h0e9d: o_data_a = 16'b1110001100001000;
            14'h0e9e: o_data_a = 16'b0000000000000011;
            14'h0e9f: o_data_a = 16'b1111110111100000;
            14'h0ea0: o_data_a = 16'b1110110111100000;
            14'h0ea1: o_data_a = 16'b1111110000010000;
            14'h0ea2: o_data_a = 16'b0000000000000000;
            14'h0ea3: o_data_a = 16'b1111110111101000;
            14'h0ea4: o_data_a = 16'b1110110010100000;
            14'h0ea5: o_data_a = 16'b1110001100001000;
            14'h0ea6: o_data_a = 16'b0000000000000000;
            14'h0ea7: o_data_a = 16'b1111110010101000;
            14'h0ea8: o_data_a = 16'b1111110000010000;
            14'h0ea9: o_data_a = 16'b1110110010100000;
            14'h0eaa: o_data_a = 16'b1111000010001000;
            14'h0eab: o_data_a = 16'b0000000000000011;
            14'h0eac: o_data_a = 16'b1110110000010000;
            14'h0ead: o_data_a = 16'b0000000000000000;
            14'h0eae: o_data_a = 16'b1111110111101000;
            14'h0eaf: o_data_a = 16'b1110110010100000;
            14'h0eb0: o_data_a = 16'b1110001100001000;
            14'h0eb1: o_data_a = 16'b0000000000000000;
            14'h0eb2: o_data_a = 16'b1111110010101000;
            14'h0eb3: o_data_a = 16'b1111110000010000;
            14'h0eb4: o_data_a = 16'b1110110010100000;
            14'h0eb5: o_data_a = 16'b1111000111001000;
            14'h0eb6: o_data_a = 16'b0000000000000011;
            14'h0eb7: o_data_a = 16'b1111110111100000;
            14'h0eb8: o_data_a = 16'b1111110000010000;
            14'h0eb9: o_data_a = 16'b0000000000000000;
            14'h0eba: o_data_a = 16'b1111110111101000;
            14'h0ebb: o_data_a = 16'b1110110010100000;
            14'h0ebc: o_data_a = 16'b1110001100001000;
            14'h0ebd: o_data_a = 16'b0000000000000011;
            14'h0ebe: o_data_a = 16'b1111110000100000;
            14'h0ebf: o_data_a = 16'b1111110000010000;
            14'h0ec0: o_data_a = 16'b0000000000000000;
            14'h0ec1: o_data_a = 16'b1111110111101000;
            14'h0ec2: o_data_a = 16'b1110110010100000;
            14'h0ec3: o_data_a = 16'b1110001100001000;
            14'h0ec4: o_data_a = 16'b0000000000000011;
            14'h0ec5: o_data_a = 16'b1111110111100000;
            14'h0ec6: o_data_a = 16'b1110110111100000;
            14'h0ec7: o_data_a = 16'b1111110000010000;
            14'h0ec8: o_data_a = 16'b0000000000000000;
            14'h0ec9: o_data_a = 16'b1111110111101000;
            14'h0eca: o_data_a = 16'b1110110010100000;
            14'h0ecb: o_data_a = 16'b1110001100001000;
            14'h0ecc: o_data_a = 16'b0000000000000000;
            14'h0ecd: o_data_a = 16'b1111110010101000;
            14'h0ece: o_data_a = 16'b1111110000010000;
            14'h0ecf: o_data_a = 16'b1110110010100000;
            14'h0ed0: o_data_a = 16'b1111000010001000;
            14'h0ed1: o_data_a = 16'b0000000000000011;
            14'h0ed2: o_data_a = 16'b1111110111100000;
            14'h0ed3: o_data_a = 16'b1111110000010000;
            14'h0ed4: o_data_a = 16'b0000000000000000;
            14'h0ed5: o_data_a = 16'b1111110111101000;
            14'h0ed6: o_data_a = 16'b1110110010100000;
            14'h0ed7: o_data_a = 16'b1110001100001000;
            14'h0ed8: o_data_a = 16'b0000000000000011;
            14'h0ed9: o_data_a = 16'b1111110000010000;
            14'h0eda: o_data_a = 16'b0000000000000011;
            14'h0edb: o_data_a = 16'b1110000010100000;
            14'h0edc: o_data_a = 16'b1111110000010000;
            14'h0edd: o_data_a = 16'b0000000000000000;
            14'h0ede: o_data_a = 16'b1111110111101000;
            14'h0edf: o_data_a = 16'b1110110010100000;
            14'h0ee0: o_data_a = 16'b1110001100001000;
            14'h0ee1: o_data_a = 16'b0000000000000000;
            14'h0ee2: o_data_a = 16'b1111110010101000;
            14'h0ee3: o_data_a = 16'b1111110000010000;
            14'h0ee4: o_data_a = 16'b1110110010100000;
            14'h0ee5: o_data_a = 16'b1111000010001000;
            14'h0ee6: o_data_a = 16'b0000000000000100;
            14'h0ee7: o_data_a = 16'b1110110000010000;
            14'h0ee8: o_data_a = 16'b0000000000001101;
            14'h0ee9: o_data_a = 16'b1110001100001000;
            14'h0eea: o_data_a = 16'b0101011101010010;
            14'h0eeb: o_data_a = 16'b1110110000010000;
            14'h0eec: o_data_a = 16'b0000000000001110;
            14'h0eed: o_data_a = 16'b1110001100001000;
            14'h0eee: o_data_a = 16'b0000111011110010;
            14'h0eef: o_data_a = 16'b1110110000010000;
            14'h0ef0: o_data_a = 16'b0000000001011111;
            14'h0ef1: o_data_a = 16'b1110101010000111;
            14'h0ef2: o_data_a = 16'b0000000000000000;
            14'h0ef3: o_data_a = 16'b1111110010101000;
            14'h0ef4: o_data_a = 16'b1111110000010000;
            14'h0ef5: o_data_a = 16'b0000000000000101;
            14'h0ef6: o_data_a = 16'b1110001100001000;
            14'h0ef7: o_data_a = 16'b0000000000000000;
            14'h0ef8: o_data_a = 16'b1111110111001000;
            14'h0ef9: o_data_a = 16'b1111110010100000;
            14'h0efa: o_data_a = 16'b1110101010001000;
            14'h0efb: o_data_a = 16'b0000000000110110;
            14'h0efc: o_data_a = 16'b1110101010000111;
            14'h0efd: o_data_a = 16'b0000000000000000;
            14'h0efe: o_data_a = 16'b1111110111101000;
            14'h0eff: o_data_a = 16'b1110110010100000;
            14'h0f00: o_data_a = 16'b1110101010001000;
            14'h0f01: o_data_a = 16'b0000000000000000;
            14'h0f02: o_data_a = 16'b1110110000010000;
            14'h0f03: o_data_a = 16'b0000000000001101;
            14'h0f04: o_data_a = 16'b1110001100001000;
            14'h0f05: o_data_a = 16'b0001000110011100;
            14'h0f06: o_data_a = 16'b1110110000010000;
            14'h0f07: o_data_a = 16'b0000000000001110;
            14'h0f08: o_data_a = 16'b1110001100001000;
            14'h0f09: o_data_a = 16'b0000111100001101;
            14'h0f0a: o_data_a = 16'b1110110000010000;
            14'h0f0b: o_data_a = 16'b0000000001011111;
            14'h0f0c: o_data_a = 16'b1110101010000111;
            14'h0f0d: o_data_a = 16'b0000000000000000;
            14'h0f0e: o_data_a = 16'b1111110010101000;
            14'h0f0f: o_data_a = 16'b1111110000010000;
            14'h0f10: o_data_a = 16'b0000000000000101;
            14'h0f11: o_data_a = 16'b1110001100001000;
            14'h0f12: o_data_a = 16'b0000000000000000;
            14'h0f13: o_data_a = 16'b1110110000010000;
            14'h0f14: o_data_a = 16'b0000000000001101;
            14'h0f15: o_data_a = 16'b1110001100001000;
            14'h0f16: o_data_a = 16'b0001000110110011;
            14'h0f17: o_data_a = 16'b1110110000010000;
            14'h0f18: o_data_a = 16'b0000000000001110;
            14'h0f19: o_data_a = 16'b1110001100001000;
            14'h0f1a: o_data_a = 16'b0000111100011110;
            14'h0f1b: o_data_a = 16'b1110110000010000;
            14'h0f1c: o_data_a = 16'b0000000001011111;
            14'h0f1d: o_data_a = 16'b1110101010000111;
            14'h0f1e: o_data_a = 16'b0000000000000000;
            14'h0f1f: o_data_a = 16'b1111110010101000;
            14'h0f20: o_data_a = 16'b1111110000010000;
            14'h0f21: o_data_a = 16'b0000000000000001;
            14'h0f22: o_data_a = 16'b1111110000100000;
            14'h0f23: o_data_a = 16'b1110001100001000;
            14'h0f24: o_data_a = 16'b0000000000000001;
            14'h0f25: o_data_a = 16'b1111110000100000;
            14'h0f26: o_data_a = 16'b1111110000010000;
            14'h0f27: o_data_a = 16'b0000000000000000;
            14'h0f28: o_data_a = 16'b1111110111101000;
            14'h0f29: o_data_a = 16'b1110110010100000;
            14'h0f2a: o_data_a = 16'b1110001100001000;
            14'h0f2b: o_data_a = 16'b0000000000000001;
            14'h0f2c: o_data_a = 16'b1110110000010000;
            14'h0f2d: o_data_a = 16'b0000000000001101;
            14'h0f2e: o_data_a = 16'b1110001100001000;
            14'h0f2f: o_data_a = 16'b0001000110111011;
            14'h0f30: o_data_a = 16'b1110110000010000;
            14'h0f31: o_data_a = 16'b0000000000001110;
            14'h0f32: o_data_a = 16'b1110001100001000;
            14'h0f33: o_data_a = 16'b0000111100110111;
            14'h0f34: o_data_a = 16'b1110110000010000;
            14'h0f35: o_data_a = 16'b0000000001011111;
            14'h0f36: o_data_a = 16'b1110101010000111;
            14'h0f37: o_data_a = 16'b0000000000000000;
            14'h0f38: o_data_a = 16'b1111110010101000;
            14'h0f39: o_data_a = 16'b1111110000010000;
            14'h0f3a: o_data_a = 16'b0000000000000101;
            14'h0f3b: o_data_a = 16'b1110001100001000;
            14'h0f3c: o_data_a = 16'b0000000000000001;
            14'h0f3d: o_data_a = 16'b1111110000100000;
            14'h0f3e: o_data_a = 16'b1111110000010000;
            14'h0f3f: o_data_a = 16'b0000000000000000;
            14'h0f40: o_data_a = 16'b1111110111101000;
            14'h0f41: o_data_a = 16'b1110110010100000;
            14'h0f42: o_data_a = 16'b1110001100001000;
            14'h0f43: o_data_a = 16'b0000000000000001;
            14'h0f44: o_data_a = 16'b1110110000010000;
            14'h0f45: o_data_a = 16'b0000000000001101;
            14'h0f46: o_data_a = 16'b1110001100001000;
            14'h0f47: o_data_a = 16'b0001000101000011;
            14'h0f48: o_data_a = 16'b1110110000010000;
            14'h0f49: o_data_a = 16'b0000000000001110;
            14'h0f4a: o_data_a = 16'b1110001100001000;
            14'h0f4b: o_data_a = 16'b0000111101001111;
            14'h0f4c: o_data_a = 16'b1110110000010000;
            14'h0f4d: o_data_a = 16'b0000000001011111;
            14'h0f4e: o_data_a = 16'b1110101010000111;
            14'h0f4f: o_data_a = 16'b0000000000000000;
            14'h0f50: o_data_a = 16'b1111110010101000;
            14'h0f51: o_data_a = 16'b1111110000010000;
            14'h0f52: o_data_a = 16'b0000000000000101;
            14'h0f53: o_data_a = 16'b1110001100001000;
            14'h0f54: o_data_a = 16'b0000000000000000;
            14'h0f55: o_data_a = 16'b1111110111001000;
            14'h0f56: o_data_a = 16'b1111110010100000;
            14'h0f57: o_data_a = 16'b1110101010001000;
            14'h0f58: o_data_a = 16'b0000000000110110;
            14'h0f59: o_data_a = 16'b1110101010000111;
            14'h0f5a: o_data_a = 16'b0000000000000111;
            14'h0f5b: o_data_a = 16'b1110110000010000;
            14'h0f5c: o_data_a = 16'b0000000000000000;
            14'h0f5d: o_data_a = 16'b1111110111101000;
            14'h0f5e: o_data_a = 16'b1110110010100000;
            14'h0f5f: o_data_a = 16'b1110001100001000;
            14'h0f60: o_data_a = 16'b0000000000000001;
            14'h0f61: o_data_a = 16'b1110110000010000;
            14'h0f62: o_data_a = 16'b0000000000001101;
            14'h0f63: o_data_a = 16'b1110001100001000;
            14'h0f64: o_data_a = 16'b0010000111000011;
            14'h0f65: o_data_a = 16'b1110110000010000;
            14'h0f66: o_data_a = 16'b0000000000001110;
            14'h0f67: o_data_a = 16'b1110001100001000;
            14'h0f68: o_data_a = 16'b0000111101101100;
            14'h0f69: o_data_a = 16'b1110110000010000;
            14'h0f6a: o_data_a = 16'b0000000001011111;
            14'h0f6b: o_data_a = 16'b1110101010000111;
            14'h0f6c: o_data_a = 16'b0000000000000000;
            14'h0f6d: o_data_a = 16'b1111110010101000;
            14'h0f6e: o_data_a = 16'b1111110000010000;
            14'h0f6f: o_data_a = 16'b0000000000000011;
            14'h0f70: o_data_a = 16'b1110001100001000;
            14'h0f71: o_data_a = 16'b0000000000000000;
            14'h0f72: o_data_a = 16'b1110110000010000;
            14'h0f73: o_data_a = 16'b0000000000001101;
            14'h0f74: o_data_a = 16'b1110001100001000;
            14'h0f75: o_data_a = 16'b0101000001110110;
            14'h0f76: o_data_a = 16'b1110110000010000;
            14'h0f77: o_data_a = 16'b0000000000001110;
            14'h0f78: o_data_a = 16'b1110001100001000;
            14'h0f79: o_data_a = 16'b0000111101111101;
            14'h0f7a: o_data_a = 16'b1110110000010000;
            14'h0f7b: o_data_a = 16'b0000000001011111;
            14'h0f7c: o_data_a = 16'b1110101010000111;
            14'h0f7d: o_data_a = 16'b0000000000000000;
            14'h0f7e: o_data_a = 16'b1111110010101000;
            14'h0f7f: o_data_a = 16'b1111110000010000;
            14'h0f80: o_data_a = 16'b0000000000000101;
            14'h0f81: o_data_a = 16'b1110001100001000;
            14'h0f82: o_data_a = 16'b0000000000110010;
            14'h0f83: o_data_a = 16'b1110110000010000;
            14'h0f84: o_data_a = 16'b0000000000000000;
            14'h0f85: o_data_a = 16'b1111110111101000;
            14'h0f86: o_data_a = 16'b1110110010100000;
            14'h0f87: o_data_a = 16'b1110001100001000;
            14'h0f88: o_data_a = 16'b0000000000000000;
            14'h0f89: o_data_a = 16'b1111110010101000;
            14'h0f8a: o_data_a = 16'b1111110000010000;
            14'h0f8b: o_data_a = 16'b0000000000000011;
            14'h0f8c: o_data_a = 16'b1111110111100000;
            14'h0f8d: o_data_a = 16'b1110110111100000;
            14'h0f8e: o_data_a = 16'b1110110111100000;
            14'h0f8f: o_data_a = 16'b1110110111100000;
            14'h0f90: o_data_a = 16'b1110110111100000;
            14'h0f91: o_data_a = 16'b1110110111100000;
            14'h0f92: o_data_a = 16'b1110001100001000;
            14'h0f93: o_data_a = 16'b0000000011100110;
            14'h0f94: o_data_a = 16'b1110110000010000;
            14'h0f95: o_data_a = 16'b0000000000000000;
            14'h0f96: o_data_a = 16'b1111110111101000;
            14'h0f97: o_data_a = 16'b1110110010100000;
            14'h0f98: o_data_a = 16'b1110001100001000;
            14'h0f99: o_data_a = 16'b0000000011100101;
            14'h0f9a: o_data_a = 16'b1110110000010000;
            14'h0f9b: o_data_a = 16'b0000000000000000;
            14'h0f9c: o_data_a = 16'b1111110111101000;
            14'h0f9d: o_data_a = 16'b1110110010100000;
            14'h0f9e: o_data_a = 16'b1110001100001000;
            14'h0f9f: o_data_a = 16'b0000000000000011;
            14'h0fa0: o_data_a = 16'b1111110000010000;
            14'h0fa1: o_data_a = 16'b0000000000000110;
            14'h0fa2: o_data_a = 16'b1110000010100000;
            14'h0fa3: o_data_a = 16'b1111110000010000;
            14'h0fa4: o_data_a = 16'b0000000000000000;
            14'h0fa5: o_data_a = 16'b1111110111101000;
            14'h0fa6: o_data_a = 16'b1110110010100000;
            14'h0fa7: o_data_a = 16'b1110001100001000;
            14'h0fa8: o_data_a = 16'b0000000000000111;
            14'h0fa9: o_data_a = 16'b1110110000010000;
            14'h0faa: o_data_a = 16'b0000000000000000;
            14'h0fab: o_data_a = 16'b1111110111101000;
            14'h0fac: o_data_a = 16'b1110110010100000;
            14'h0fad: o_data_a = 16'b1110001100001000;
            14'h0fae: o_data_a = 16'b0000000000000100;
            14'h0faf: o_data_a = 16'b1110110000010000;
            14'h0fb0: o_data_a = 16'b0000000000001101;
            14'h0fb1: o_data_a = 16'b1110001100001000;
            14'h0fb2: o_data_a = 16'b0000101001100011;
            14'h0fb3: o_data_a = 16'b1110110000010000;
            14'h0fb4: o_data_a = 16'b0000000000001110;
            14'h0fb5: o_data_a = 16'b1110001100001000;
            14'h0fb6: o_data_a = 16'b0000111110111010;
            14'h0fb7: o_data_a = 16'b1110110000010000;
            14'h0fb8: o_data_a = 16'b0000000001011111;
            14'h0fb9: o_data_a = 16'b1110101010000111;
            14'h0fba: o_data_a = 16'b0000000000000000;
            14'h0fbb: o_data_a = 16'b1111110010101000;
            14'h0fbc: o_data_a = 16'b1111110000010000;
            14'h0fbd: o_data_a = 16'b0000000000000011;
            14'h0fbe: o_data_a = 16'b1111110000100000;
            14'h0fbf: o_data_a = 16'b1110001100001000;
            14'h0fc0: o_data_a = 16'b0000000011111101;
            14'h0fc1: o_data_a = 16'b1110110000010000;
            14'h0fc2: o_data_a = 16'b0000000000000000;
            14'h0fc3: o_data_a = 16'b1111110111101000;
            14'h0fc4: o_data_a = 16'b1110110010100000;
            14'h0fc5: o_data_a = 16'b1110001100001000;
            14'h0fc6: o_data_a = 16'b0000000011011110;
            14'h0fc7: o_data_a = 16'b1110110000010000;
            14'h0fc8: o_data_a = 16'b0000000000000000;
            14'h0fc9: o_data_a = 16'b1111110111101000;
            14'h0fca: o_data_a = 16'b1110110010100000;
            14'h0fcb: o_data_a = 16'b1110001100001000;
            14'h0fcc: o_data_a = 16'b0000000000000000;
            14'h0fcd: o_data_a = 16'b1111110111001000;
            14'h0fce: o_data_a = 16'b1111110010100000;
            14'h0fcf: o_data_a = 16'b1110101010001000;
            14'h0fd0: o_data_a = 16'b0000000111111111;
            14'h0fd1: o_data_a = 16'b1110110000010000;
            14'h0fd2: o_data_a = 16'b0000000000000000;
            14'h0fd3: o_data_a = 16'b1111110111101000;
            14'h0fd4: o_data_a = 16'b1110110010100000;
            14'h0fd5: o_data_a = 16'b1110001100001000;
            14'h0fd6: o_data_a = 16'b0000000000000000;
            14'h0fd7: o_data_a = 16'b1111110111001000;
            14'h0fd8: o_data_a = 16'b1111110010100000;
            14'h0fd9: o_data_a = 16'b1110101010001000;
            14'h0fda: o_data_a = 16'b0000000011100101;
            14'h0fdb: o_data_a = 16'b1110110000010000;
            14'h0fdc: o_data_a = 16'b0000000000000000;
            14'h0fdd: o_data_a = 16'b1111110111101000;
            14'h0fde: o_data_a = 16'b1110110010100000;
            14'h0fdf: o_data_a = 16'b1110001100001000;
            14'h0fe0: o_data_a = 16'b0000000000000110;
            14'h0fe1: o_data_a = 16'b1110110000010000;
            14'h0fe2: o_data_a = 16'b0000000000001101;
            14'h0fe3: o_data_a = 16'b1110001100001000;
            14'h0fe4: o_data_a = 16'b0000000010010001;
            14'h0fe5: o_data_a = 16'b1110110000010000;
            14'h0fe6: o_data_a = 16'b0000000000001110;
            14'h0fe7: o_data_a = 16'b1110001100001000;
            14'h0fe8: o_data_a = 16'b0000111111101100;
            14'h0fe9: o_data_a = 16'b1110110000010000;
            14'h0fea: o_data_a = 16'b0000000001011111;
            14'h0feb: o_data_a = 16'b1110101010000111;
            14'h0fec: o_data_a = 16'b0000000000000000;
            14'h0fed: o_data_a = 16'b1111110010101000;
            14'h0fee: o_data_a = 16'b1111110000010000;
            14'h0fef: o_data_a = 16'b0000000000000011;
            14'h0ff0: o_data_a = 16'b1111110111100000;
            14'h0ff1: o_data_a = 16'b1110001100001000;
            14'h0ff2: o_data_a = 16'b0000000000000011;
            14'h0ff3: o_data_a = 16'b1111110111100000;
            14'h0ff4: o_data_a = 16'b1111110000010000;
            14'h0ff5: o_data_a = 16'b0000000000000000;
            14'h0ff6: o_data_a = 16'b1111110111101000;
            14'h0ff7: o_data_a = 16'b1110110010100000;
            14'h0ff8: o_data_a = 16'b1110001100001000;
            14'h0ff9: o_data_a = 16'b0000000110010000;
            14'h0ffa: o_data_a = 16'b1110110000010000;
            14'h0ffb: o_data_a = 16'b0000000000000000;
            14'h0ffc: o_data_a = 16'b1111110111101000;
            14'h0ffd: o_data_a = 16'b1110110010100000;
            14'h0ffe: o_data_a = 16'b1110001100001000;
            14'h0fff: o_data_a = 16'b0000000000000000;
            14'h1000: o_data_a = 16'b1111110111001000;
            14'h1001: o_data_a = 16'b1111110010100000;
            14'h1002: o_data_a = 16'b1110101010001000;
            14'h1003: o_data_a = 16'b0000000000000011;
            14'h1004: o_data_a = 16'b1110110000010000;
            14'h1005: o_data_a = 16'b0000000000001101;
            14'h1006: o_data_a = 16'b1110001100001000;
            14'h1007: o_data_a = 16'b0000001010001100;
            14'h1008: o_data_a = 16'b1110110000010000;
            14'h1009: o_data_a = 16'b0000000000001110;
            14'h100a: o_data_a = 16'b1110001100001000;
            14'h100b: o_data_a = 16'b0001000000001111;
            14'h100c: o_data_a = 16'b1110110000010000;
            14'h100d: o_data_a = 16'b0000000001011111;
            14'h100e: o_data_a = 16'b1110101010000111;
            14'h100f: o_data_a = 16'b0000000000000000;
            14'h1010: o_data_a = 16'b1111110010101000;
            14'h1011: o_data_a = 16'b1111110000010000;
            14'h1012: o_data_a = 16'b0000000000000101;
            14'h1013: o_data_a = 16'b1110001100001000;
            14'h1014: o_data_a = 16'b0000000000000000;
            14'h1015: o_data_a = 16'b1111110111001000;
            14'h1016: o_data_a = 16'b1111110010100000;
            14'h1017: o_data_a = 16'b1110101010001000;
            14'h1018: o_data_a = 16'b0000000011101110;
            14'h1019: o_data_a = 16'b1110110000010000;
            14'h101a: o_data_a = 16'b0000000000000000;
            14'h101b: o_data_a = 16'b1111110111101000;
            14'h101c: o_data_a = 16'b1110110010100000;
            14'h101d: o_data_a = 16'b1110001100001000;
            14'h101e: o_data_a = 16'b0000000111111111;
            14'h101f: o_data_a = 16'b1110110000010000;
            14'h1020: o_data_a = 16'b0000000000000000;
            14'h1021: o_data_a = 16'b1111110111101000;
            14'h1022: o_data_a = 16'b1110110010100000;
            14'h1023: o_data_a = 16'b1110001100001000;
            14'h1024: o_data_a = 16'b0000000011110000;
            14'h1025: o_data_a = 16'b1110110000010000;
            14'h1026: o_data_a = 16'b0000000000000000;
            14'h1027: o_data_a = 16'b1111110111101000;
            14'h1028: o_data_a = 16'b1110110010100000;
            14'h1029: o_data_a = 16'b1110001100001000;
            14'h102a: o_data_a = 16'b0000000000000100;
            14'h102b: o_data_a = 16'b1110110000010000;
            14'h102c: o_data_a = 16'b0000000000001101;
            14'h102d: o_data_a = 16'b1110001100001000;
            14'h102e: o_data_a = 16'b0101011101010010;
            14'h102f: o_data_a = 16'b1110110000010000;
            14'h1030: o_data_a = 16'b0000000000001110;
            14'h1031: o_data_a = 16'b1110001100001000;
            14'h1032: o_data_a = 16'b0001000000110110;
            14'h1033: o_data_a = 16'b1110110000010000;
            14'h1034: o_data_a = 16'b0000000001011111;
            14'h1035: o_data_a = 16'b1110101010000111;
            14'h1036: o_data_a = 16'b0000000000000000;
            14'h1037: o_data_a = 16'b1111110010101000;
            14'h1038: o_data_a = 16'b1111110000010000;
            14'h1039: o_data_a = 16'b0000000000000101;
            14'h103a: o_data_a = 16'b1110001100001000;
            14'h103b: o_data_a = 16'b0000000000010110;
            14'h103c: o_data_a = 16'b1110110000010000;
            14'h103d: o_data_a = 16'b0000000000000000;
            14'h103e: o_data_a = 16'b1111110111101000;
            14'h103f: o_data_a = 16'b1110110010100000;
            14'h1040: o_data_a = 16'b1110001100001000;
            14'h1041: o_data_a = 16'b0000000000000000;
            14'h1042: o_data_a = 16'b1111110111001000;
            14'h1043: o_data_a = 16'b1111110010100000;
            14'h1044: o_data_a = 16'b1110101010001000;
            14'h1045: o_data_a = 16'b0000000000000010;
            14'h1046: o_data_a = 16'b1110110000010000;
            14'h1047: o_data_a = 16'b0000000000001101;
            14'h1048: o_data_a = 16'b1110001100001000;
            14'h1049: o_data_a = 16'b0100101110010110;
            14'h104a: o_data_a = 16'b1110110000010000;
            14'h104b: o_data_a = 16'b0000000000001110;
            14'h104c: o_data_a = 16'b1110001100001000;
            14'h104d: o_data_a = 16'b0001000001010001;
            14'h104e: o_data_a = 16'b1110110000010000;
            14'h104f: o_data_a = 16'b0000000001011111;
            14'h1050: o_data_a = 16'b1110101010000111;
            14'h1051: o_data_a = 16'b0000000000000000;
            14'h1052: o_data_a = 16'b1111110010101000;
            14'h1053: o_data_a = 16'b1111110000010000;
            14'h1054: o_data_a = 16'b0000000000000101;
            14'h1055: o_data_a = 16'b1110001100001000;
            14'h1056: o_data_a = 16'b0000000000001000;
            14'h1057: o_data_a = 16'b1110110000010000;
            14'h1058: o_data_a = 16'b0000000000000000;
            14'h1059: o_data_a = 16'b1111110111101000;
            14'h105a: o_data_a = 16'b1110110010100000;
            14'h105b: o_data_a = 16'b1110001100001000;
            14'h105c: o_data_a = 16'b0000000000000001;
            14'h105d: o_data_a = 16'b1110110000010000;
            14'h105e: o_data_a = 16'b0000000000001101;
            14'h105f: o_data_a = 16'b1110001100001000;
            14'h1060: o_data_a = 16'b0110001000010001;
            14'h1061: o_data_a = 16'b1110110000010000;
            14'h1062: o_data_a = 16'b0000000000001110;
            14'h1063: o_data_a = 16'b1110001100001000;
            14'h1064: o_data_a = 16'b0001000001101000;
            14'h1065: o_data_a = 16'b1110110000010000;
            14'h1066: o_data_a = 16'b0000000001011111;
            14'h1067: o_data_a = 16'b1110101010000111;
            14'h1068: o_data_a = 16'b0000000001010011;
            14'h1069: o_data_a = 16'b1110110000010000;
            14'h106a: o_data_a = 16'b0000000000000000;
            14'h106b: o_data_a = 16'b1111110111101000;
            14'h106c: o_data_a = 16'b1110110010100000;
            14'h106d: o_data_a = 16'b1110001100001000;
            14'h106e: o_data_a = 16'b0000000000000010;
            14'h106f: o_data_a = 16'b1110110000010000;
            14'h1070: o_data_a = 16'b0000000000001101;
            14'h1071: o_data_a = 16'b1110001100001000;
            14'h1072: o_data_a = 16'b0110010000111011;
            14'h1073: o_data_a = 16'b1110110000010000;
            14'h1074: o_data_a = 16'b0000000000001110;
            14'h1075: o_data_a = 16'b1110001100001000;
            14'h1076: o_data_a = 16'b0001000001111010;
            14'h1077: o_data_a = 16'b1110110000010000;
            14'h1078: o_data_a = 16'b0000000001011111;
            14'h1079: o_data_a = 16'b1110101010000111;
            14'h107a: o_data_a = 16'b0000000001100011;
            14'h107b: o_data_a = 16'b1110110000010000;
            14'h107c: o_data_a = 16'b0000000000000000;
            14'h107d: o_data_a = 16'b1111110111101000;
            14'h107e: o_data_a = 16'b1110110010100000;
            14'h107f: o_data_a = 16'b1110001100001000;
            14'h1080: o_data_a = 16'b0000000000000010;
            14'h1081: o_data_a = 16'b1110110000010000;
            14'h1082: o_data_a = 16'b0000000000001101;
            14'h1083: o_data_a = 16'b1110001100001000;
            14'h1084: o_data_a = 16'b0110010000111011;
            14'h1085: o_data_a = 16'b1110110000010000;
            14'h1086: o_data_a = 16'b0000000000001110;
            14'h1087: o_data_a = 16'b1110001100001000;
            14'h1088: o_data_a = 16'b0001000010001100;
            14'h1089: o_data_a = 16'b1110110000010000;
            14'h108a: o_data_a = 16'b0000000001011111;
            14'h108b: o_data_a = 16'b1110101010000111;
            14'h108c: o_data_a = 16'b0000000001101111;
            14'h108d: o_data_a = 16'b1110110000010000;
            14'h108e: o_data_a = 16'b0000000000000000;
            14'h108f: o_data_a = 16'b1111110111101000;
            14'h1090: o_data_a = 16'b1110110010100000;
            14'h1091: o_data_a = 16'b1110001100001000;
            14'h1092: o_data_a = 16'b0000000000000010;
            14'h1093: o_data_a = 16'b1110110000010000;
            14'h1094: o_data_a = 16'b0000000000001101;
            14'h1095: o_data_a = 16'b1110001100001000;
            14'h1096: o_data_a = 16'b0110010000111011;
            14'h1097: o_data_a = 16'b1110110000010000;
            14'h1098: o_data_a = 16'b0000000000001110;
            14'h1099: o_data_a = 16'b1110001100001000;
            14'h109a: o_data_a = 16'b0001000010011110;
            14'h109b: o_data_a = 16'b1110110000010000;
            14'h109c: o_data_a = 16'b0000000001011111;
            14'h109d: o_data_a = 16'b1110101010000111;
            14'h109e: o_data_a = 16'b0000000001110010;
            14'h109f: o_data_a = 16'b1110110000010000;
            14'h10a0: o_data_a = 16'b0000000000000000;
            14'h10a1: o_data_a = 16'b1111110111101000;
            14'h10a2: o_data_a = 16'b1110110010100000;
            14'h10a3: o_data_a = 16'b1110001100001000;
            14'h10a4: o_data_a = 16'b0000000000000010;
            14'h10a5: o_data_a = 16'b1110110000010000;
            14'h10a6: o_data_a = 16'b0000000000001101;
            14'h10a7: o_data_a = 16'b1110001100001000;
            14'h10a8: o_data_a = 16'b0110010000111011;
            14'h10a9: o_data_a = 16'b1110110000010000;
            14'h10aa: o_data_a = 16'b0000000000001110;
            14'h10ab: o_data_a = 16'b1110001100001000;
            14'h10ac: o_data_a = 16'b0001000010110000;
            14'h10ad: o_data_a = 16'b1110110000010000;
            14'h10ae: o_data_a = 16'b0000000001011111;
            14'h10af: o_data_a = 16'b1110101010000111;
            14'h10b0: o_data_a = 16'b0000000001100101;
            14'h10b1: o_data_a = 16'b1110110000010000;
            14'h10b2: o_data_a = 16'b0000000000000000;
            14'h10b3: o_data_a = 16'b1111110111101000;
            14'h10b4: o_data_a = 16'b1110110010100000;
            14'h10b5: o_data_a = 16'b1110001100001000;
            14'h10b6: o_data_a = 16'b0000000000000010;
            14'h10b7: o_data_a = 16'b1110110000010000;
            14'h10b8: o_data_a = 16'b0000000000001101;
            14'h10b9: o_data_a = 16'b1110001100001000;
            14'h10ba: o_data_a = 16'b0110010000111011;
            14'h10bb: o_data_a = 16'b1110110000010000;
            14'h10bc: o_data_a = 16'b0000000000001110;
            14'h10bd: o_data_a = 16'b1110001100001000;
            14'h10be: o_data_a = 16'b0001000011000010;
            14'h10bf: o_data_a = 16'b1110110000010000;
            14'h10c0: o_data_a = 16'b0000000001011111;
            14'h10c1: o_data_a = 16'b1110101010000111;
            14'h10c2: o_data_a = 16'b0000000000111010;
            14'h10c3: o_data_a = 16'b1110110000010000;
            14'h10c4: o_data_a = 16'b0000000000000000;
            14'h10c5: o_data_a = 16'b1111110111101000;
            14'h10c6: o_data_a = 16'b1110110010100000;
            14'h10c7: o_data_a = 16'b1110001100001000;
            14'h10c8: o_data_a = 16'b0000000000000010;
            14'h10c9: o_data_a = 16'b1110110000010000;
            14'h10ca: o_data_a = 16'b0000000000001101;
            14'h10cb: o_data_a = 16'b1110001100001000;
            14'h10cc: o_data_a = 16'b0110010000111011;
            14'h10cd: o_data_a = 16'b1110110000010000;
            14'h10ce: o_data_a = 16'b0000000000001110;
            14'h10cf: o_data_a = 16'b1110001100001000;
            14'h10d0: o_data_a = 16'b0001000011010100;
            14'h10d1: o_data_a = 16'b1110110000010000;
            14'h10d2: o_data_a = 16'b0000000001011111;
            14'h10d3: o_data_a = 16'b1110101010000111;
            14'h10d4: o_data_a = 16'b0000000000100000;
            14'h10d5: o_data_a = 16'b1110110000010000;
            14'h10d6: o_data_a = 16'b0000000000000000;
            14'h10d7: o_data_a = 16'b1111110111101000;
            14'h10d8: o_data_a = 16'b1110110010100000;
            14'h10d9: o_data_a = 16'b1110001100001000;
            14'h10da: o_data_a = 16'b0000000000000010;
            14'h10db: o_data_a = 16'b1110110000010000;
            14'h10dc: o_data_a = 16'b0000000000001101;
            14'h10dd: o_data_a = 16'b1110001100001000;
            14'h10de: o_data_a = 16'b0110010000111011;
            14'h10df: o_data_a = 16'b1110110000010000;
            14'h10e0: o_data_a = 16'b0000000000001110;
            14'h10e1: o_data_a = 16'b1110001100001000;
            14'h10e2: o_data_a = 16'b0001000011100110;
            14'h10e3: o_data_a = 16'b1110110000010000;
            14'h10e4: o_data_a = 16'b0000000001011111;
            14'h10e5: o_data_a = 16'b1110101010000111;
            14'h10e6: o_data_a = 16'b0000000000110000;
            14'h10e7: o_data_a = 16'b1110110000010000;
            14'h10e8: o_data_a = 16'b0000000000000000;
            14'h10e9: o_data_a = 16'b1111110111101000;
            14'h10ea: o_data_a = 16'b1110110010100000;
            14'h10eb: o_data_a = 16'b1110001100001000;
            14'h10ec: o_data_a = 16'b0000000000000010;
            14'h10ed: o_data_a = 16'b1110110000010000;
            14'h10ee: o_data_a = 16'b0000000000001101;
            14'h10ef: o_data_a = 16'b1110001100001000;
            14'h10f0: o_data_a = 16'b0110010000111011;
            14'h10f1: o_data_a = 16'b1110110000010000;
            14'h10f2: o_data_a = 16'b0000000000001110;
            14'h10f3: o_data_a = 16'b1110001100001000;
            14'h10f4: o_data_a = 16'b0001000011111000;
            14'h10f5: o_data_a = 16'b1110110000010000;
            14'h10f6: o_data_a = 16'b0000000001011111;
            14'h10f7: o_data_a = 16'b1110101010000111;
            14'h10f8: o_data_a = 16'b0000000000000001;
            14'h10f9: o_data_a = 16'b1110110000010000;
            14'h10fa: o_data_a = 16'b0000000000001101;
            14'h10fb: o_data_a = 16'b1110001100001000;
            14'h10fc: o_data_a = 16'b0100110110001010;
            14'h10fd: o_data_a = 16'b1110110000010000;
            14'h10fe: o_data_a = 16'b0000000000001110;
            14'h10ff: o_data_a = 16'b1110001100001000;
            14'h1100: o_data_a = 16'b0001000100000100;
            14'h1101: o_data_a = 16'b1110110000010000;
            14'h1102: o_data_a = 16'b0000000001011111;
            14'h1103: o_data_a = 16'b1110101010000111;
            14'h1104: o_data_a = 16'b0000000000000000;
            14'h1105: o_data_a = 16'b1111110010101000;
            14'h1106: o_data_a = 16'b1111110000010000;
            14'h1107: o_data_a = 16'b0000000000000101;
            14'h1108: o_data_a = 16'b1110001100001000;
            14'h1109: o_data_a = 16'b0000000000000000;
            14'h110a: o_data_a = 16'b1111110111001000;
            14'h110b: o_data_a = 16'b1111110010100000;
            14'h110c: o_data_a = 16'b1110101010001000;
            14'h110d: o_data_a = 16'b0000000000000000;
            14'h110e: o_data_a = 16'b1111110010101000;
            14'h110f: o_data_a = 16'b1111110000010000;
            14'h1110: o_data_a = 16'b0000000000000011;
            14'h1111: o_data_a = 16'b1111110111100000;
            14'h1112: o_data_a = 16'b1110110111100000;
            14'h1113: o_data_a = 16'b1110110111100000;
            14'h1114: o_data_a = 16'b1110001100001000;
            14'h1115: o_data_a = 16'b0000000000000000;
            14'h1116: o_data_a = 16'b1111110111001000;
            14'h1117: o_data_a = 16'b1111110010100000;
            14'h1118: o_data_a = 16'b1110101010001000;
            14'h1119: o_data_a = 16'b0000000000000000;
            14'h111a: o_data_a = 16'b1111110010101000;
            14'h111b: o_data_a = 16'b1111110000010000;
            14'h111c: o_data_a = 16'b0000000000000011;
            14'h111d: o_data_a = 16'b1111110111100000;
            14'h111e: o_data_a = 16'b1110110111100000;
            14'h111f: o_data_a = 16'b1110110111100000;
            14'h1120: o_data_a = 16'b1110110111100000;
            14'h1121: o_data_a = 16'b1110001100001000;
            14'h1122: o_data_a = 16'b0000000000000000;
            14'h1123: o_data_a = 16'b1111110111001000;
            14'h1124: o_data_a = 16'b1111110010100000;
            14'h1125: o_data_a = 16'b1110101010001000;
            14'h1126: o_data_a = 16'b0000000000000000;
            14'h1127: o_data_a = 16'b1111110010101000;
            14'h1128: o_data_a = 16'b1111110000010000;
            14'h1129: o_data_a = 16'b0000000000000011;
            14'h112a: o_data_a = 16'b1111110111100000;
            14'h112b: o_data_a = 16'b1110110111100000;
            14'h112c: o_data_a = 16'b1110001100001000;
            14'h112d: o_data_a = 16'b0000000000000000;
            14'h112e: o_data_a = 16'b1111110111001000;
            14'h112f: o_data_a = 16'b1111110010100000;
            14'h1130: o_data_a = 16'b1110101010001000;
            14'h1131: o_data_a = 16'b0000000000000000;
            14'h1132: o_data_a = 16'b1111110010101000;
            14'h1133: o_data_a = 16'b1111110000010000;
            14'h1134: o_data_a = 16'b0000000000000011;
            14'h1135: o_data_a = 16'b1111110111100000;
            14'h1136: o_data_a = 16'b1110110111100000;
            14'h1137: o_data_a = 16'b1110110111100000;
            14'h1138: o_data_a = 16'b1110110111100000;
            14'h1139: o_data_a = 16'b1110110111100000;
            14'h113a: o_data_a = 16'b1110001100001000;
            14'h113b: o_data_a = 16'b0000000000000011;
            14'h113c: o_data_a = 16'b1111110000010000;
            14'h113d: o_data_a = 16'b0000000000000000;
            14'h113e: o_data_a = 16'b1111110111101000;
            14'h113f: o_data_a = 16'b1110110010100000;
            14'h1140: o_data_a = 16'b1110001100001000;
            14'h1141: o_data_a = 16'b0000000000110110;
            14'h1142: o_data_a = 16'b1110101010000111;
            14'h1143: o_data_a = 16'b0000000000000010;
            14'h1144: o_data_a = 16'b1111110000100000;
            14'h1145: o_data_a = 16'b1111110000010000;
            14'h1146: o_data_a = 16'b0000000000000000;
            14'h1147: o_data_a = 16'b1111110111101000;
            14'h1148: o_data_a = 16'b1110110010100000;
            14'h1149: o_data_a = 16'b1110001100001000;
            14'h114a: o_data_a = 16'b0000000000000000;
            14'h114b: o_data_a = 16'b1111110010101000;
            14'h114c: o_data_a = 16'b1111110000010000;
            14'h114d: o_data_a = 16'b0000000000000011;
            14'h114e: o_data_a = 16'b1110001100001000;
            14'h114f: o_data_a = 16'b0000000000000011;
            14'h1150: o_data_a = 16'b1111110000100000;
            14'h1151: o_data_a = 16'b1111110000010000;
            14'h1152: o_data_a = 16'b0000000000000000;
            14'h1153: o_data_a = 16'b1111110111101000;
            14'h1154: o_data_a = 16'b1110110010100000;
            14'h1155: o_data_a = 16'b1110001100001000;
            14'h1156: o_data_a = 16'b0000000000000001;
            14'h1157: o_data_a = 16'b1110110000010000;
            14'h1158: o_data_a = 16'b0000000000001101;
            14'h1159: o_data_a = 16'b1110001100001000;
            14'h115a: o_data_a = 16'b0000101011100010;
            14'h115b: o_data_a = 16'b1110110000010000;
            14'h115c: o_data_a = 16'b0000000000001110;
            14'h115d: o_data_a = 16'b1110001100001000;
            14'h115e: o_data_a = 16'b0001000101100010;
            14'h115f: o_data_a = 16'b1110110000010000;
            14'h1160: o_data_a = 16'b0000000001011111;
            14'h1161: o_data_a = 16'b1110101010000111;
            14'h1162: o_data_a = 16'b0000000000000000;
            14'h1163: o_data_a = 16'b1111110010101000;
            14'h1164: o_data_a = 16'b1111110000010000;
            14'h1165: o_data_a = 16'b0000000000000101;
            14'h1166: o_data_a = 16'b1110001100001000;
            14'h1167: o_data_a = 16'b0000000000000011;
            14'h1168: o_data_a = 16'b1111110111100000;
            14'h1169: o_data_a = 16'b1111110000010000;
            14'h116a: o_data_a = 16'b0000000000000000;
            14'h116b: o_data_a = 16'b1111110111101000;
            14'h116c: o_data_a = 16'b1110110010100000;
            14'h116d: o_data_a = 16'b1110001100001000;
            14'h116e: o_data_a = 16'b0000000000000001;
            14'h116f: o_data_a = 16'b1110110000010000;
            14'h1170: o_data_a = 16'b0000000000001101;
            14'h1171: o_data_a = 16'b1110001100001000;
            14'h1172: o_data_a = 16'b0000000101011010;
            14'h1173: o_data_a = 16'b1110110000010000;
            14'h1174: o_data_a = 16'b0000000000001110;
            14'h1175: o_data_a = 16'b1110001100001000;
            14'h1176: o_data_a = 16'b0001000101111010;
            14'h1177: o_data_a = 16'b1110110000010000;
            14'h1178: o_data_a = 16'b0000000001011111;
            14'h1179: o_data_a = 16'b1110101010000111;
            14'h117a: o_data_a = 16'b0000000000000000;
            14'h117b: o_data_a = 16'b1111110010101000;
            14'h117c: o_data_a = 16'b1111110000010000;
            14'h117d: o_data_a = 16'b0000000000000101;
            14'h117e: o_data_a = 16'b1110001100001000;
            14'h117f: o_data_a = 16'b0000000000000011;
            14'h1180: o_data_a = 16'b1111110000010000;
            14'h1181: o_data_a = 16'b0000000000000000;
            14'h1182: o_data_a = 16'b1111110111101000;
            14'h1183: o_data_a = 16'b1110110010100000;
            14'h1184: o_data_a = 16'b1110001100001000;
            14'h1185: o_data_a = 16'b0000000000000001;
            14'h1186: o_data_a = 16'b1110110000010000;
            14'h1187: o_data_a = 16'b0000000000001101;
            14'h1188: o_data_a = 16'b1110001100001000;
            14'h1189: o_data_a = 16'b0010010010001101;
            14'h118a: o_data_a = 16'b1110110000010000;
            14'h118b: o_data_a = 16'b0000000000001110;
            14'h118c: o_data_a = 16'b1110001100001000;
            14'h118d: o_data_a = 16'b0001000110010001;
            14'h118e: o_data_a = 16'b1110110000010000;
            14'h118f: o_data_a = 16'b0000000001011111;
            14'h1190: o_data_a = 16'b1110101010000111;
            14'h1191: o_data_a = 16'b0000000000000000;
            14'h1192: o_data_a = 16'b1111110010101000;
            14'h1193: o_data_a = 16'b1111110000010000;
            14'h1194: o_data_a = 16'b0000000000000101;
            14'h1195: o_data_a = 16'b1110001100001000;
            14'h1196: o_data_a = 16'b0000000000000000;
            14'h1197: o_data_a = 16'b1111110111001000;
            14'h1198: o_data_a = 16'b1111110010100000;
            14'h1199: o_data_a = 16'b1110101010001000;
            14'h119a: o_data_a = 16'b0000000000110110;
            14'h119b: o_data_a = 16'b1110101010000111;
            14'h119c: o_data_a = 16'b0000000000000000;
            14'h119d: o_data_a = 16'b1110110000010000;
            14'h119e: o_data_a = 16'b0000000000001101;
            14'h119f: o_data_a = 16'b1110001100001000;
            14'h11a0: o_data_a = 16'b0000111101011010;
            14'h11a1: o_data_a = 16'b1110110000010000;
            14'h11a2: o_data_a = 16'b0000000000001110;
            14'h11a3: o_data_a = 16'b1110001100001000;
            14'h11a4: o_data_a = 16'b0001000110101000;
            14'h11a5: o_data_a = 16'b1110110000010000;
            14'h11a6: o_data_a = 16'b0000000001011111;
            14'h11a7: o_data_a = 16'b1110101010000111;
            14'h11a8: o_data_a = 16'b0000000000000000;
            14'h11a9: o_data_a = 16'b1111110010101000;
            14'h11aa: o_data_a = 16'b1111110000010000;
            14'h11ab: o_data_a = 16'b0000000000010000;
            14'h11ac: o_data_a = 16'b1110001100001000;
            14'h11ad: o_data_a = 16'b0000000000000000;
            14'h11ae: o_data_a = 16'b1111110111001000;
            14'h11af: o_data_a = 16'b1111110010100000;
            14'h11b0: o_data_a = 16'b1110101010001000;
            14'h11b1: o_data_a = 16'b0000000000110110;
            14'h11b2: o_data_a = 16'b1110101010000111;
            14'h11b3: o_data_a = 16'b0000000000010000;
            14'h11b4: o_data_a = 16'b1111110000010000;
            14'h11b5: o_data_a = 16'b0000000000000000;
            14'h11b6: o_data_a = 16'b1111110111101000;
            14'h11b7: o_data_a = 16'b1110110010100000;
            14'h11b8: o_data_a = 16'b1110001100001000;
            14'h11b9: o_data_a = 16'b0000000000110110;
            14'h11ba: o_data_a = 16'b1110101010000111;
            14'h11bb: o_data_a = 16'b0000000000000000;
            14'h11bc: o_data_a = 16'b1111110111101000;
            14'h11bd: o_data_a = 16'b1110110010100000;
            14'h11be: o_data_a = 16'b1110101010001000;
            14'h11bf: o_data_a = 16'b0000000000000010;
            14'h11c0: o_data_a = 16'b1111110000100000;
            14'h11c1: o_data_a = 16'b1111110000010000;
            14'h11c2: o_data_a = 16'b0000000000000000;
            14'h11c3: o_data_a = 16'b1111110111101000;
            14'h11c4: o_data_a = 16'b1110110010100000;
            14'h11c5: o_data_a = 16'b1110001100001000;
            14'h11c6: o_data_a = 16'b0000000000000000;
            14'h11c7: o_data_a = 16'b1111110010101000;
            14'h11c8: o_data_a = 16'b1111110000010000;
            14'h11c9: o_data_a = 16'b0000000000000011;
            14'h11ca: o_data_a = 16'b1110001100001000;
            14'h11cb: o_data_a = 16'b0000000000000011;
            14'h11cc: o_data_a = 16'b1111110000010000;
            14'h11cd: o_data_a = 16'b0000000000000011;
            14'h11ce: o_data_a = 16'b1110000010100000;
            14'h11cf: o_data_a = 16'b1111110000010000;
            14'h11d0: o_data_a = 16'b0000000000000000;
            14'h11d1: o_data_a = 16'b1111110111101000;
            14'h11d2: o_data_a = 16'b1110110010100000;
            14'h11d3: o_data_a = 16'b1110001100001000;
            14'h11d4: o_data_a = 16'b0000000000000000;
            14'h11d5: o_data_a = 16'b1111110010100000;
            14'h11d6: o_data_a = 16'b1111110001001000;
            14'h11d7: o_data_a = 16'b0000000000000000;
            14'h11d8: o_data_a = 16'b1111110010100000;
            14'h11d9: o_data_a = 16'b1111110001001000;
            14'h11da: o_data_a = 16'b0000000000000000;
            14'h11db: o_data_a = 16'b1111110010101000;
            14'h11dc: o_data_a = 16'b1111110000010000;
            14'h11dd: o_data_a = 16'b0001001101001111;
            14'h11de: o_data_a = 16'b1110001100000101;
            14'h11df: o_data_a = 16'b0000000000000001;
            14'h11e0: o_data_a = 16'b1111110000100000;
            14'h11e1: o_data_a = 16'b1111110000010000;
            14'h11e2: o_data_a = 16'b0000000000000000;
            14'h11e3: o_data_a = 16'b1111110111101000;
            14'h11e4: o_data_a = 16'b1110110010100000;
            14'h11e5: o_data_a = 16'b1110001100001000;
            14'h11e6: o_data_a = 16'b0000000000000000;
            14'h11e7: o_data_a = 16'b1111110111001000;
            14'h11e8: o_data_a = 16'b1111110010100000;
            14'h11e9: o_data_a = 16'b1110101010001000;
            14'h11ea: o_data_a = 16'b0001000111101110;
            14'h11eb: o_data_a = 16'b1110110000010000;
            14'h11ec: o_data_a = 16'b0000000000000110;
            14'h11ed: o_data_a = 16'b1110101010000111;
            14'h11ee: o_data_a = 16'b0000000000000011;
            14'h11ef: o_data_a = 16'b1111110000010000;
            14'h11f0: o_data_a = 16'b0000000000000011;
            14'h11f1: o_data_a = 16'b1110000010100000;
            14'h11f2: o_data_a = 16'b1111110000010000;
            14'h11f3: o_data_a = 16'b0000000000000000;
            14'h11f4: o_data_a = 16'b1111110111101000;
            14'h11f5: o_data_a = 16'b1110110010100000;
            14'h11f6: o_data_a = 16'b1110001100001000;
            14'h11f7: o_data_a = 16'b0000000000000000;
            14'h11f8: o_data_a = 16'b1111110010100000;
            14'h11f9: o_data_a = 16'b1111110001001000;
            14'h11fa: o_data_a = 16'b0000000000000000;
            14'h11fb: o_data_a = 16'b1111110010101000;
            14'h11fc: o_data_a = 16'b1111110000010000;
            14'h11fd: o_data_a = 16'b1110110010100000;
            14'h11fe: o_data_a = 16'b1111000000001000;
            14'h11ff: o_data_a = 16'b0000000000000000;
            14'h1200: o_data_a = 16'b1111110010100000;
            14'h1201: o_data_a = 16'b1111110001001000;
            14'h1202: o_data_a = 16'b0000000000000000;
            14'h1203: o_data_a = 16'b1111110010101000;
            14'h1204: o_data_a = 16'b1111110000010000;
            14'h1205: o_data_a = 16'b0001001001001010;
            14'h1206: o_data_a = 16'b1110001100000101;
            14'h1207: o_data_a = 16'b0000000000000000;
            14'h1208: o_data_a = 16'b1110110000010000;
            14'h1209: o_data_a = 16'b0000000000001101;
            14'h120a: o_data_a = 16'b1110001100001000;
            14'h120b: o_data_a = 16'b0001011100100100;
            14'h120c: o_data_a = 16'b1110110000010000;
            14'h120d: o_data_a = 16'b0000000000001110;
            14'h120e: o_data_a = 16'b1110001100001000;
            14'h120f: o_data_a = 16'b0001001000010011;
            14'h1210: o_data_a = 16'b1110110000010000;
            14'h1211: o_data_a = 16'b0000000001011111;
            14'h1212: o_data_a = 16'b1110101010000111;
            14'h1213: o_data_a = 16'b0000000000000000;
            14'h1214: o_data_a = 16'b1111110010101000;
            14'h1215: o_data_a = 16'b1111110000010000;
            14'h1216: o_data_a = 16'b0000000000000001;
            14'h1217: o_data_a = 16'b1111110000100000;
            14'h1218: o_data_a = 16'b1110001100001000;
            14'h1219: o_data_a = 16'b0000000000000011;
            14'h121a: o_data_a = 16'b1111110000100000;
            14'h121b: o_data_a = 16'b1111110000010000;
            14'h121c: o_data_a = 16'b0000000000000000;
            14'h121d: o_data_a = 16'b1111110111101000;
            14'h121e: o_data_a = 16'b1110110010100000;
            14'h121f: o_data_a = 16'b1110001100001000;
            14'h1220: o_data_a = 16'b0000000000000001;
            14'h1221: o_data_a = 16'b1110110000010000;
            14'h1222: o_data_a = 16'b0000000000001101;
            14'h1223: o_data_a = 16'b1110001100001000;
            14'h1224: o_data_a = 16'b0000110010001011;
            14'h1225: o_data_a = 16'b1110110000010000;
            14'h1226: o_data_a = 16'b0000000000001110;
            14'h1227: o_data_a = 16'b1110001100001000;
            14'h1228: o_data_a = 16'b0001001000101100;
            14'h1229: o_data_a = 16'b1110110000010000;
            14'h122a: o_data_a = 16'b0000000001011111;
            14'h122b: o_data_a = 16'b1110101010000111;
            14'h122c: o_data_a = 16'b0000000000000000;
            14'h122d: o_data_a = 16'b1111110010101000;
            14'h122e: o_data_a = 16'b1111110000010000;
            14'h122f: o_data_a = 16'b0000000000000101;
            14'h1230: o_data_a = 16'b1110001100001000;
            14'h1231: o_data_a = 16'b0000000000000011;
            14'h1232: o_data_a = 16'b1111110000010000;
            14'h1233: o_data_a = 16'b0000000000000000;
            14'h1234: o_data_a = 16'b1111110111101000;
            14'h1235: o_data_a = 16'b1110110010100000;
            14'h1236: o_data_a = 16'b1110001100001000;
            14'h1237: o_data_a = 16'b0000000000000001;
            14'h1238: o_data_a = 16'b1110110000010000;
            14'h1239: o_data_a = 16'b0000000000001101;
            14'h123a: o_data_a = 16'b1110001100001000;
            14'h123b: o_data_a = 16'b0001010001000111;
            14'h123c: o_data_a = 16'b1110110000010000;
            14'h123d: o_data_a = 16'b0000000000001110;
            14'h123e: o_data_a = 16'b1110001100001000;
            14'h123f: o_data_a = 16'b0001001001000011;
            14'h1240: o_data_a = 16'b1110110000010000;
            14'h1241: o_data_a = 16'b0000000001011111;
            14'h1242: o_data_a = 16'b1110101010000111;
            14'h1243: o_data_a = 16'b0000000000000000;
            14'h1244: o_data_a = 16'b1111110010101000;
            14'h1245: o_data_a = 16'b1111110000010000;
            14'h1246: o_data_a = 16'b0000000000000101;
            14'h1247: o_data_a = 16'b1110001100001000;
            14'h1248: o_data_a = 16'b0001000111011111;
            14'h1249: o_data_a = 16'b1110101010000111;
            14'h124a: o_data_a = 16'b0000000000000001;
            14'h124b: o_data_a = 16'b1111110000100000;
            14'h124c: o_data_a = 16'b1111110000010000;
            14'h124d: o_data_a = 16'b0000000000000000;
            14'h124e: o_data_a = 16'b1111110111101000;
            14'h124f: o_data_a = 16'b1110110010100000;
            14'h1250: o_data_a = 16'b1110001100001000;
            14'h1251: o_data_a = 16'b0000000010000010;
            14'h1252: o_data_a = 16'b1110110000010000;
            14'h1253: o_data_a = 16'b0000000000000000;
            14'h1254: o_data_a = 16'b1111110111101000;
            14'h1255: o_data_a = 16'b1110110010100000;
            14'h1256: o_data_a = 16'b1110001100001000;
            14'h1257: o_data_a = 16'b0001001001011011;
            14'h1258: o_data_a = 16'b1110110000010000;
            14'h1259: o_data_a = 16'b0000000000000110;
            14'h125a: o_data_a = 16'b1110101010000111;
            14'h125b: o_data_a = 16'b0000000000000000;
            14'h125c: o_data_a = 16'b1111110010101000;
            14'h125d: o_data_a = 16'b1111110000010000;
            14'h125e: o_data_a = 16'b0001001001100010;
            14'h125f: o_data_a = 16'b1110001100000101;
            14'h1260: o_data_a = 16'b0001001010000000;
            14'h1261: o_data_a = 16'b1110101010000111;
            14'h1262: o_data_a = 16'b0000000000000011;
            14'h1263: o_data_a = 16'b1111110000100000;
            14'h1264: o_data_a = 16'b1111110000010000;
            14'h1265: o_data_a = 16'b0000000000000000;
            14'h1266: o_data_a = 16'b1111110111101000;
            14'h1267: o_data_a = 16'b1110110010100000;
            14'h1268: o_data_a = 16'b1110001100001000;
            14'h1269: o_data_a = 16'b0000000000000000;
            14'h126a: o_data_a = 16'b1111110111001000;
            14'h126b: o_data_a = 16'b1111110010100000;
            14'h126c: o_data_a = 16'b1110111111001000;
            14'h126d: o_data_a = 16'b0000000000000010;
            14'h126e: o_data_a = 16'b1110110000010000;
            14'h126f: o_data_a = 16'b0000000000001101;
            14'h1270: o_data_a = 16'b1110001100001000;
            14'h1271: o_data_a = 16'b0000101111100100;
            14'h1272: o_data_a = 16'b1110110000010000;
            14'h1273: o_data_a = 16'b0000000000001110;
            14'h1274: o_data_a = 16'b1110001100001000;
            14'h1275: o_data_a = 16'b0001001001111001;
            14'h1276: o_data_a = 16'b1110110000010000;
            14'h1277: o_data_a = 16'b0000000001011111;
            14'h1278: o_data_a = 16'b1110101010000111;
            14'h1279: o_data_a = 16'b0000000000000000;
            14'h127a: o_data_a = 16'b1111110010101000;
            14'h127b: o_data_a = 16'b1111110000010000;
            14'h127c: o_data_a = 16'b0000000000000101;
            14'h127d: o_data_a = 16'b1110001100001000;
            14'h127e: o_data_a = 16'b0001001011011111;
            14'h127f: o_data_a = 16'b1110101010000111;
            14'h1280: o_data_a = 16'b0000000000000001;
            14'h1281: o_data_a = 16'b1111110000100000;
            14'h1282: o_data_a = 16'b1111110000010000;
            14'h1283: o_data_a = 16'b0000000000000000;
            14'h1284: o_data_a = 16'b1111110111101000;
            14'h1285: o_data_a = 16'b1110110010100000;
            14'h1286: o_data_a = 16'b1110001100001000;
            14'h1287: o_data_a = 16'b0000000010000100;
            14'h1288: o_data_a = 16'b1110110000010000;
            14'h1289: o_data_a = 16'b0000000000000000;
            14'h128a: o_data_a = 16'b1111110111101000;
            14'h128b: o_data_a = 16'b1110110010100000;
            14'h128c: o_data_a = 16'b1110001100001000;
            14'h128d: o_data_a = 16'b0001001010010001;
            14'h128e: o_data_a = 16'b1110110000010000;
            14'h128f: o_data_a = 16'b0000000000000110;
            14'h1290: o_data_a = 16'b1110101010000111;
            14'h1291: o_data_a = 16'b0000000000000000;
            14'h1292: o_data_a = 16'b1111110010101000;
            14'h1293: o_data_a = 16'b1111110000010000;
            14'h1294: o_data_a = 16'b0001001010011000;
            14'h1295: o_data_a = 16'b1110001100000101;
            14'h1296: o_data_a = 16'b0001001010111000;
            14'h1297: o_data_a = 16'b1110101010000111;
            14'h1298: o_data_a = 16'b0000000000000011;
            14'h1299: o_data_a = 16'b1111110000100000;
            14'h129a: o_data_a = 16'b1111110000010000;
            14'h129b: o_data_a = 16'b0000000000000000;
            14'h129c: o_data_a = 16'b1111110111101000;
            14'h129d: o_data_a = 16'b1110110010100000;
            14'h129e: o_data_a = 16'b1110001100001000;
            14'h129f: o_data_a = 16'b0000000000000010;
            14'h12a0: o_data_a = 16'b1110110000010000;
            14'h12a1: o_data_a = 16'b0000000000000000;
            14'h12a2: o_data_a = 16'b1111110111101000;
            14'h12a3: o_data_a = 16'b1110110010100000;
            14'h12a4: o_data_a = 16'b1110001100001000;
            14'h12a5: o_data_a = 16'b0000000000000010;
            14'h12a6: o_data_a = 16'b1110110000010000;
            14'h12a7: o_data_a = 16'b0000000000001101;
            14'h12a8: o_data_a = 16'b1110001100001000;
            14'h12a9: o_data_a = 16'b0000101111100100;
            14'h12aa: o_data_a = 16'b1110110000010000;
            14'h12ab: o_data_a = 16'b0000000000001110;
            14'h12ac: o_data_a = 16'b1110001100001000;
            14'h12ad: o_data_a = 16'b0001001010110001;
            14'h12ae: o_data_a = 16'b1110110000010000;
            14'h12af: o_data_a = 16'b0000000001011111;
            14'h12b0: o_data_a = 16'b1110101010000111;
            14'h12b1: o_data_a = 16'b0000000000000000;
            14'h12b2: o_data_a = 16'b1111110010101000;
            14'h12b3: o_data_a = 16'b1111110000010000;
            14'h12b4: o_data_a = 16'b0000000000000101;
            14'h12b5: o_data_a = 16'b1110001100001000;
            14'h12b6: o_data_a = 16'b0001001011011111;
            14'h12b7: o_data_a = 16'b1110101010000111;
            14'h12b8: o_data_a = 16'b0000000000000001;
            14'h12b9: o_data_a = 16'b1111110000100000;
            14'h12ba: o_data_a = 16'b1111110000010000;
            14'h12bb: o_data_a = 16'b0000000000000000;
            14'h12bc: o_data_a = 16'b1111110111101000;
            14'h12bd: o_data_a = 16'b1110110010100000;
            14'h12be: o_data_a = 16'b1110001100001000;
            14'h12bf: o_data_a = 16'b0000000010001100;
            14'h12c0: o_data_a = 16'b1110110000010000;
            14'h12c1: o_data_a = 16'b0000000000000000;
            14'h12c2: o_data_a = 16'b1111110111101000;
            14'h12c3: o_data_a = 16'b1110110010100000;
            14'h12c4: o_data_a = 16'b1110001100001000;
            14'h12c5: o_data_a = 16'b0001001011001001;
            14'h12c6: o_data_a = 16'b1110110000010000;
            14'h12c7: o_data_a = 16'b0000000000000110;
            14'h12c8: o_data_a = 16'b1110101010000111;
            14'h12c9: o_data_a = 16'b0000000000000000;
            14'h12ca: o_data_a = 16'b1111110010101000;
            14'h12cb: o_data_a = 16'b1111110000010000;
            14'h12cc: o_data_a = 16'b0001001011010000;
            14'h12cd: o_data_a = 16'b1110001100000101;
            14'h12ce: o_data_a = 16'b0001001011011111;
            14'h12cf: o_data_a = 16'b1110101010000111;
            14'h12d0: o_data_a = 16'b0000000000000000;
            14'h12d1: o_data_a = 16'b1111110111001000;
            14'h12d2: o_data_a = 16'b1111110010100000;
            14'h12d3: o_data_a = 16'b1110101010001000;
            14'h12d4: o_data_a = 16'b0000000000000000;
            14'h12d5: o_data_a = 16'b1111110010100000;
            14'h12d6: o_data_a = 16'b1111110001001000;
            14'h12d7: o_data_a = 16'b0000000000000000;
            14'h12d8: o_data_a = 16'b1111110010101000;
            14'h12d9: o_data_a = 16'b1111110000010000;
            14'h12da: o_data_a = 16'b0000000000000011;
            14'h12db: o_data_a = 16'b1111110111100000;
            14'h12dc: o_data_a = 16'b1110110111100000;
            14'h12dd: o_data_a = 16'b1110110111100000;
            14'h12de: o_data_a = 16'b1110001100001000;
            14'h12df: o_data_a = 16'b0000000000000001;
            14'h12e0: o_data_a = 16'b1111110000100000;
            14'h12e1: o_data_a = 16'b1111110000010000;
            14'h12e2: o_data_a = 16'b0000000000000000;
            14'h12e3: o_data_a = 16'b1111110111101000;
            14'h12e4: o_data_a = 16'b1110110010100000;
            14'h12e5: o_data_a = 16'b1110001100001000;
            14'h12e6: o_data_a = 16'b0000000000000000;
            14'h12e7: o_data_a = 16'b1111110111001000;
            14'h12e8: o_data_a = 16'b1111110010100000;
            14'h12e9: o_data_a = 16'b1110101010001000;
            14'h12ea: o_data_a = 16'b0001001011101110;
            14'h12eb: o_data_a = 16'b1110110000010000;
            14'h12ec: o_data_a = 16'b0000000000000110;
            14'h12ed: o_data_a = 16'b1110101010000111;
            14'h12ee: o_data_a = 16'b0000000000000000;
            14'h12ef: o_data_a = 16'b1111110010100000;
            14'h12f0: o_data_a = 16'b1111110001001000;
            14'h12f1: o_data_a = 16'b0000000000000011;
            14'h12f2: o_data_a = 16'b1111110000010000;
            14'h12f3: o_data_a = 16'b0000000000000011;
            14'h12f4: o_data_a = 16'b1110000010100000;
            14'h12f5: o_data_a = 16'b1111110000010000;
            14'h12f6: o_data_a = 16'b0000000000000000;
            14'h12f7: o_data_a = 16'b1111110111101000;
            14'h12f8: o_data_a = 16'b1110110010100000;
            14'h12f9: o_data_a = 16'b1110001100001000;
            14'h12fa: o_data_a = 16'b0000000000000000;
            14'h12fb: o_data_a = 16'b1111110010100000;
            14'h12fc: o_data_a = 16'b1111110001001000;
            14'h12fd: o_data_a = 16'b0000000000000000;
            14'h12fe: o_data_a = 16'b1111110010101000;
            14'h12ff: o_data_a = 16'b1111110000010000;
            14'h1300: o_data_a = 16'b1110110010100000;
            14'h1301: o_data_a = 16'b1111000000001000;
            14'h1302: o_data_a = 16'b0000000000000000;
            14'h1303: o_data_a = 16'b1111110010100000;
            14'h1304: o_data_a = 16'b1111110001001000;
            14'h1305: o_data_a = 16'b0000000000000000;
            14'h1306: o_data_a = 16'b1111110010101000;
            14'h1307: o_data_a = 16'b1111110000010000;
            14'h1308: o_data_a = 16'b0001001101001101;
            14'h1309: o_data_a = 16'b1110001100000101;
            14'h130a: o_data_a = 16'b0000000000000000;
            14'h130b: o_data_a = 16'b1110110000010000;
            14'h130c: o_data_a = 16'b0000000000001101;
            14'h130d: o_data_a = 16'b1110001100001000;
            14'h130e: o_data_a = 16'b0001011100100100;
            14'h130f: o_data_a = 16'b1110110000010000;
            14'h1310: o_data_a = 16'b0000000000001110;
            14'h1311: o_data_a = 16'b1110001100001000;
            14'h1312: o_data_a = 16'b0001001100010110;
            14'h1313: o_data_a = 16'b1110110000010000;
            14'h1314: o_data_a = 16'b0000000001011111;
            14'h1315: o_data_a = 16'b1110101010000111;
            14'h1316: o_data_a = 16'b0000000000000000;
            14'h1317: o_data_a = 16'b1111110010101000;
            14'h1318: o_data_a = 16'b1111110000010000;
            14'h1319: o_data_a = 16'b0000000000000001;
            14'h131a: o_data_a = 16'b1111110000100000;
            14'h131b: o_data_a = 16'b1110001100001000;
            14'h131c: o_data_a = 16'b0000000000000011;
            14'h131d: o_data_a = 16'b1111110000100000;
            14'h131e: o_data_a = 16'b1111110000010000;
            14'h131f: o_data_a = 16'b0000000000000000;
            14'h1320: o_data_a = 16'b1111110111101000;
            14'h1321: o_data_a = 16'b1110110010100000;
            14'h1322: o_data_a = 16'b1110001100001000;
            14'h1323: o_data_a = 16'b0000000000000001;
            14'h1324: o_data_a = 16'b1110110000010000;
            14'h1325: o_data_a = 16'b0000000000001101;
            14'h1326: o_data_a = 16'b1110001100001000;
            14'h1327: o_data_a = 16'b0000110010001011;
            14'h1328: o_data_a = 16'b1110110000010000;
            14'h1329: o_data_a = 16'b0000000000001110;
            14'h132a: o_data_a = 16'b1110001100001000;
            14'h132b: o_data_a = 16'b0001001100101111;
            14'h132c: o_data_a = 16'b1110110000010000;
            14'h132d: o_data_a = 16'b0000000001011111;
            14'h132e: o_data_a = 16'b1110101010000111;
            14'h132f: o_data_a = 16'b0000000000000000;
            14'h1330: o_data_a = 16'b1111110010101000;
            14'h1331: o_data_a = 16'b1111110000010000;
            14'h1332: o_data_a = 16'b0000000000000101;
            14'h1333: o_data_a = 16'b1110001100001000;
            14'h1334: o_data_a = 16'b0000000000000011;
            14'h1335: o_data_a = 16'b1111110000010000;
            14'h1336: o_data_a = 16'b0000000000000000;
            14'h1337: o_data_a = 16'b1111110111101000;
            14'h1338: o_data_a = 16'b1110110010100000;
            14'h1339: o_data_a = 16'b1110001100001000;
            14'h133a: o_data_a = 16'b0000000000000001;
            14'h133b: o_data_a = 16'b1110110000010000;
            14'h133c: o_data_a = 16'b0000000000001101;
            14'h133d: o_data_a = 16'b1110001100001000;
            14'h133e: o_data_a = 16'b0001010001000111;
            14'h133f: o_data_a = 16'b1110110000010000;
            14'h1340: o_data_a = 16'b0000000000001110;
            14'h1341: o_data_a = 16'b1110001100001000;
            14'h1342: o_data_a = 16'b0001001101000110;
            14'h1343: o_data_a = 16'b1110110000010000;
            14'h1344: o_data_a = 16'b0000000001011111;
            14'h1345: o_data_a = 16'b1110101010000111;
            14'h1346: o_data_a = 16'b0000000000000000;
            14'h1347: o_data_a = 16'b1111110010101000;
            14'h1348: o_data_a = 16'b1111110000010000;
            14'h1349: o_data_a = 16'b0000000000000101;
            14'h134a: o_data_a = 16'b1110001100001000;
            14'h134b: o_data_a = 16'b0001001011011111;
            14'h134c: o_data_a = 16'b1110101010000111;
            14'h134d: o_data_a = 16'b0001000111001011;
            14'h134e: o_data_a = 16'b1110101010000111;
            14'h134f: o_data_a = 16'b0000000000000011;
            14'h1350: o_data_a = 16'b1111110000010000;
            14'h1351: o_data_a = 16'b0000000000000011;
            14'h1352: o_data_a = 16'b1110000010100000;
            14'h1353: o_data_a = 16'b1111110000010000;
            14'h1354: o_data_a = 16'b0000000000000000;
            14'h1355: o_data_a = 16'b1111110111101000;
            14'h1356: o_data_a = 16'b1110110010100000;
            14'h1357: o_data_a = 16'b1110001100001000;
            14'h1358: o_data_a = 16'b0000000000000000;
            14'h1359: o_data_a = 16'b1111110010101000;
            14'h135a: o_data_a = 16'b1111110000010000;
            14'h135b: o_data_a = 16'b0001001101011111;
            14'h135c: o_data_a = 16'b1110001100000101;
            14'h135d: o_data_a = 16'b0001010001000001;
            14'h135e: o_data_a = 16'b1110101010000111;
            14'h135f: o_data_a = 16'b0000000000001010;
            14'h1360: o_data_a = 16'b1110110000010000;
            14'h1361: o_data_a = 16'b0000000000000000;
            14'h1362: o_data_a = 16'b1111110111101000;
            14'h1363: o_data_a = 16'b1110110010100000;
            14'h1364: o_data_a = 16'b1110001100001000;
            14'h1365: o_data_a = 16'b0000000000011011;
            14'h1366: o_data_a = 16'b1110110000010000;
            14'h1367: o_data_a = 16'b0000000000000000;
            14'h1368: o_data_a = 16'b1111110111101000;
            14'h1369: o_data_a = 16'b1110110010100000;
            14'h136a: o_data_a = 16'b1110001100001000;
            14'h136b: o_data_a = 16'b0000000000000010;
            14'h136c: o_data_a = 16'b1110110000010000;
            14'h136d: o_data_a = 16'b0000000000001101;
            14'h136e: o_data_a = 16'b1110001100001000;
            14'h136f: o_data_a = 16'b0100101110010110;
            14'h1370: o_data_a = 16'b1110110000010000;
            14'h1371: o_data_a = 16'b0000000000001110;
            14'h1372: o_data_a = 16'b1110001100001000;
            14'h1373: o_data_a = 16'b0001001101110111;
            14'h1374: o_data_a = 16'b1110110000010000;
            14'h1375: o_data_a = 16'b0000000001011111;
            14'h1376: o_data_a = 16'b1110101010000111;
            14'h1377: o_data_a = 16'b0000000000000000;
            14'h1378: o_data_a = 16'b1111110010101000;
            14'h1379: o_data_a = 16'b1111110000010000;
            14'h137a: o_data_a = 16'b0000000000000101;
            14'h137b: o_data_a = 16'b1110001100001000;
            14'h137c: o_data_a = 16'b0000000000001001;
            14'h137d: o_data_a = 16'b1110110000010000;
            14'h137e: o_data_a = 16'b0000000000000000;
            14'h137f: o_data_a = 16'b1111110111101000;
            14'h1380: o_data_a = 16'b1110110010100000;
            14'h1381: o_data_a = 16'b1110001100001000;
            14'h1382: o_data_a = 16'b0000000000000001;
            14'h1383: o_data_a = 16'b1110110000010000;
            14'h1384: o_data_a = 16'b0000000000001101;
            14'h1385: o_data_a = 16'b1110001100001000;
            14'h1386: o_data_a = 16'b0110001000010001;
            14'h1387: o_data_a = 16'b1110110000010000;
            14'h1388: o_data_a = 16'b0000000000001110;
            14'h1389: o_data_a = 16'b1110001100001000;
            14'h138a: o_data_a = 16'b0001001110001110;
            14'h138b: o_data_a = 16'b1110110000010000;
            14'h138c: o_data_a = 16'b0000000001011111;
            14'h138d: o_data_a = 16'b1110101010000111;
            14'h138e: o_data_a = 16'b0000000001000111;
            14'h138f: o_data_a = 16'b1110110000010000;
            14'h1390: o_data_a = 16'b0000000000000000;
            14'h1391: o_data_a = 16'b1111110111101000;
            14'h1392: o_data_a = 16'b1110110010100000;
            14'h1393: o_data_a = 16'b1110001100001000;
            14'h1394: o_data_a = 16'b0000000000000010;
            14'h1395: o_data_a = 16'b1110110000010000;
            14'h1396: o_data_a = 16'b0000000000001101;
            14'h1397: o_data_a = 16'b1110001100001000;
            14'h1398: o_data_a = 16'b0110010000111011;
            14'h1399: o_data_a = 16'b1110110000010000;
            14'h139a: o_data_a = 16'b0000000000001110;
            14'h139b: o_data_a = 16'b1110001100001000;
            14'h139c: o_data_a = 16'b0001001110100000;
            14'h139d: o_data_a = 16'b1110110000010000;
            14'h139e: o_data_a = 16'b0000000001011111;
            14'h139f: o_data_a = 16'b1110101010000111;
            14'h13a0: o_data_a = 16'b0000000001100001;
            14'h13a1: o_data_a = 16'b1110110000010000;
            14'h13a2: o_data_a = 16'b0000000000000000;
            14'h13a3: o_data_a = 16'b1111110111101000;
            14'h13a4: o_data_a = 16'b1110110010100000;
            14'h13a5: o_data_a = 16'b1110001100001000;
            14'h13a6: o_data_a = 16'b0000000000000010;
            14'h13a7: o_data_a = 16'b1110110000010000;
            14'h13a8: o_data_a = 16'b0000000000001101;
            14'h13a9: o_data_a = 16'b1110001100001000;
            14'h13aa: o_data_a = 16'b0110010000111011;
            14'h13ab: o_data_a = 16'b1110110000010000;
            14'h13ac: o_data_a = 16'b0000000000001110;
            14'h13ad: o_data_a = 16'b1110001100001000;
            14'h13ae: o_data_a = 16'b0001001110110010;
            14'h13af: o_data_a = 16'b1110110000010000;
            14'h13b0: o_data_a = 16'b0000000001011111;
            14'h13b1: o_data_a = 16'b1110101010000111;
            14'h13b2: o_data_a = 16'b0000000001101101;
            14'h13b3: o_data_a = 16'b1110110000010000;
            14'h13b4: o_data_a = 16'b0000000000000000;
            14'h13b5: o_data_a = 16'b1111110111101000;
            14'h13b6: o_data_a = 16'b1110110010100000;
            14'h13b7: o_data_a = 16'b1110001100001000;
            14'h13b8: o_data_a = 16'b0000000000000010;
            14'h13b9: o_data_a = 16'b1110110000010000;
            14'h13ba: o_data_a = 16'b0000000000001101;
            14'h13bb: o_data_a = 16'b1110001100001000;
            14'h13bc: o_data_a = 16'b0110010000111011;
            14'h13bd: o_data_a = 16'b1110110000010000;
            14'h13be: o_data_a = 16'b0000000000001110;
            14'h13bf: o_data_a = 16'b1110001100001000;
            14'h13c0: o_data_a = 16'b0001001111000100;
            14'h13c1: o_data_a = 16'b1110110000010000;
            14'h13c2: o_data_a = 16'b0000000001011111;
            14'h13c3: o_data_a = 16'b1110101010000111;
            14'h13c4: o_data_a = 16'b0000000001100101;
            14'h13c5: o_data_a = 16'b1110110000010000;
            14'h13c6: o_data_a = 16'b0000000000000000;
            14'h13c7: o_data_a = 16'b1111110111101000;
            14'h13c8: o_data_a = 16'b1110110010100000;
            14'h13c9: o_data_a = 16'b1110001100001000;
            14'h13ca: o_data_a = 16'b0000000000000010;
            14'h13cb: o_data_a = 16'b1110110000010000;
            14'h13cc: o_data_a = 16'b0000000000001101;
            14'h13cd: o_data_a = 16'b1110001100001000;
            14'h13ce: o_data_a = 16'b0110010000111011;
            14'h13cf: o_data_a = 16'b1110110000010000;
            14'h13d0: o_data_a = 16'b0000000000001110;
            14'h13d1: o_data_a = 16'b1110001100001000;
            14'h13d2: o_data_a = 16'b0001001111010110;
            14'h13d3: o_data_a = 16'b1110110000010000;
            14'h13d4: o_data_a = 16'b0000000001011111;
            14'h13d5: o_data_a = 16'b1110101010000111;
            14'h13d6: o_data_a = 16'b0000000000100000;
            14'h13d7: o_data_a = 16'b1110110000010000;
            14'h13d8: o_data_a = 16'b0000000000000000;
            14'h13d9: o_data_a = 16'b1111110111101000;
            14'h13da: o_data_a = 16'b1110110010100000;
            14'h13db: o_data_a = 16'b1110001100001000;
            14'h13dc: o_data_a = 16'b0000000000000010;
            14'h13dd: o_data_a = 16'b1110110000010000;
            14'h13de: o_data_a = 16'b0000000000001101;
            14'h13df: o_data_a = 16'b1110001100001000;
            14'h13e0: o_data_a = 16'b0110010000111011;
            14'h13e1: o_data_a = 16'b1110110000010000;
            14'h13e2: o_data_a = 16'b0000000000001110;
            14'h13e3: o_data_a = 16'b1110001100001000;
            14'h13e4: o_data_a = 16'b0001001111101000;
            14'h13e5: o_data_a = 16'b1110110000010000;
            14'h13e6: o_data_a = 16'b0000000001011111;
            14'h13e7: o_data_a = 16'b1110101010000111;
            14'h13e8: o_data_a = 16'b0000000001001111;
            14'h13e9: o_data_a = 16'b1110110000010000;
            14'h13ea: o_data_a = 16'b0000000000000000;
            14'h13eb: o_data_a = 16'b1111110111101000;
            14'h13ec: o_data_a = 16'b1110110010100000;
            14'h13ed: o_data_a = 16'b1110001100001000;
            14'h13ee: o_data_a = 16'b0000000000000010;
            14'h13ef: o_data_a = 16'b1110110000010000;
            14'h13f0: o_data_a = 16'b0000000000001101;
            14'h13f1: o_data_a = 16'b1110001100001000;
            14'h13f2: o_data_a = 16'b0110010000111011;
            14'h13f3: o_data_a = 16'b1110110000010000;
            14'h13f4: o_data_a = 16'b0000000000001110;
            14'h13f5: o_data_a = 16'b1110001100001000;
            14'h13f6: o_data_a = 16'b0001001111111010;
            14'h13f7: o_data_a = 16'b1110110000010000;
            14'h13f8: o_data_a = 16'b0000000001011111;
            14'h13f9: o_data_a = 16'b1110101010000111;
            14'h13fa: o_data_a = 16'b0000000001110110;
            14'h13fb: o_data_a = 16'b1110110000010000;
            14'h13fc: o_data_a = 16'b0000000000000000;
            14'h13fd: o_data_a = 16'b1111110111101000;
            14'h13fe: o_data_a = 16'b1110110010100000;
            14'h13ff: o_data_a = 16'b1110001100001000;
            14'h1400: o_data_a = 16'b0000000000000010;
            14'h1401: o_data_a = 16'b1110110000010000;
            14'h1402: o_data_a = 16'b0000000000001101;
            14'h1403: o_data_a = 16'b1110001100001000;
            14'h1404: o_data_a = 16'b0110010000111011;
            14'h1405: o_data_a = 16'b1110110000010000;
            14'h1406: o_data_a = 16'b0000000000001110;
            14'h1407: o_data_a = 16'b1110001100001000;
            14'h1408: o_data_a = 16'b0001010000001100;
            14'h1409: o_data_a = 16'b1110110000010000;
            14'h140a: o_data_a = 16'b0000000001011111;
            14'h140b: o_data_a = 16'b1110101010000111;
            14'h140c: o_data_a = 16'b0000000001100101;
            14'h140d: o_data_a = 16'b1110110000010000;
            14'h140e: o_data_a = 16'b0000000000000000;
            14'h140f: o_data_a = 16'b1111110111101000;
            14'h1410: o_data_a = 16'b1110110010100000;
            14'h1411: o_data_a = 16'b1110001100001000;
            14'h1412: o_data_a = 16'b0000000000000010;
            14'h1413: o_data_a = 16'b1110110000010000;
            14'h1414: o_data_a = 16'b0000000000001101;
            14'h1415: o_data_a = 16'b1110001100001000;
            14'h1416: o_data_a = 16'b0110010000111011;
            14'h1417: o_data_a = 16'b1110110000010000;
            14'h1418: o_data_a = 16'b0000000000001110;
            14'h1419: o_data_a = 16'b1110001100001000;
            14'h141a: o_data_a = 16'b0001010000011110;
            14'h141b: o_data_a = 16'b1110110000010000;
            14'h141c: o_data_a = 16'b0000000001011111;
            14'h141d: o_data_a = 16'b1110101010000111;
            14'h141e: o_data_a = 16'b0000000001110010;
            14'h141f: o_data_a = 16'b1110110000010000;
            14'h1420: o_data_a = 16'b0000000000000000;
            14'h1421: o_data_a = 16'b1111110111101000;
            14'h1422: o_data_a = 16'b1110110010100000;
            14'h1423: o_data_a = 16'b1110001100001000;
            14'h1424: o_data_a = 16'b0000000000000010;
            14'h1425: o_data_a = 16'b1110110000010000;
            14'h1426: o_data_a = 16'b0000000000001101;
            14'h1427: o_data_a = 16'b1110001100001000;
            14'h1428: o_data_a = 16'b0110010000111011;
            14'h1429: o_data_a = 16'b1110110000010000;
            14'h142a: o_data_a = 16'b0000000000001110;
            14'h142b: o_data_a = 16'b1110001100001000;
            14'h142c: o_data_a = 16'b0001010000110000;
            14'h142d: o_data_a = 16'b1110110000010000;
            14'h142e: o_data_a = 16'b0000000001011111;
            14'h142f: o_data_a = 16'b1110101010000111;
            14'h1430: o_data_a = 16'b0000000000000001;
            14'h1431: o_data_a = 16'b1110110000010000;
            14'h1432: o_data_a = 16'b0000000000001101;
            14'h1433: o_data_a = 16'b1110001100001000;
            14'h1434: o_data_a = 16'b0100110110001010;
            14'h1435: o_data_a = 16'b1110110000010000;
            14'h1436: o_data_a = 16'b0000000000001110;
            14'h1437: o_data_a = 16'b1110001100001000;
            14'h1438: o_data_a = 16'b0001010000111100;
            14'h1439: o_data_a = 16'b1110110000010000;
            14'h143a: o_data_a = 16'b0000000001011111;
            14'h143b: o_data_a = 16'b1110101010000111;
            14'h143c: o_data_a = 16'b0000000000000000;
            14'h143d: o_data_a = 16'b1111110010101000;
            14'h143e: o_data_a = 16'b1111110000010000;
            14'h143f: o_data_a = 16'b0000000000000101;
            14'h1440: o_data_a = 16'b1110001100001000;
            14'h1441: o_data_a = 16'b0000000000000000;
            14'h1442: o_data_a = 16'b1111110111001000;
            14'h1443: o_data_a = 16'b1111110010100000;
            14'h1444: o_data_a = 16'b1110101010001000;
            14'h1445: o_data_a = 16'b0000000000110110;
            14'h1446: o_data_a = 16'b1110101010000111;
            14'h1447: o_data_a = 16'b0000000000000101;
            14'h1448: o_data_a = 16'b1110110000010000;
            14'h1449: o_data_a = 16'b1110001110010000;
            14'h144a: o_data_a = 16'b0000000000000000;
            14'h144b: o_data_a = 16'b1111110111101000;
            14'h144c: o_data_a = 16'b1110110010100000;
            14'h144d: o_data_a = 16'b1110101010001000;
            14'h144e: o_data_a = 16'b0001010001001001;
            14'h144f: o_data_a = 16'b1110001100000001;
            14'h1450: o_data_a = 16'b0000000000000010;
            14'h1451: o_data_a = 16'b1111110000100000;
            14'h1452: o_data_a = 16'b1111110000010000;
            14'h1453: o_data_a = 16'b0000000000000000;
            14'h1454: o_data_a = 16'b1111110111101000;
            14'h1455: o_data_a = 16'b1110110010100000;
            14'h1456: o_data_a = 16'b1110001100001000;
            14'h1457: o_data_a = 16'b0000000000000000;
            14'h1458: o_data_a = 16'b1111110010101000;
            14'h1459: o_data_a = 16'b1111110000010000;
            14'h145a: o_data_a = 16'b0000000000000011;
            14'h145b: o_data_a = 16'b1110001100001000;
            14'h145c: o_data_a = 16'b0000000000000011;
            14'h145d: o_data_a = 16'b1111110111100000;
            14'h145e: o_data_a = 16'b1111110000010000;
            14'h145f: o_data_a = 16'b0000000000000000;
            14'h1460: o_data_a = 16'b1111110111101000;
            14'h1461: o_data_a = 16'b1110110010100000;
            14'h1462: o_data_a = 16'b1110001100001000;
            14'h1463: o_data_a = 16'b0000000000000001;
            14'h1464: o_data_a = 16'b1110110000010000;
            14'h1465: o_data_a = 16'b0000000000001101;
            14'h1466: o_data_a = 16'b1110001100001000;
            14'h1467: o_data_a = 16'b0000010001100110;
            14'h1468: o_data_a = 16'b1110110000010000;
            14'h1469: o_data_a = 16'b0000000000001110;
            14'h146a: o_data_a = 16'b1110001100001000;
            14'h146b: o_data_a = 16'b0001010001101111;
            14'h146c: o_data_a = 16'b1110110000010000;
            14'h146d: o_data_a = 16'b0000000001011111;
            14'h146e: o_data_a = 16'b1110101010000111;
            14'h146f: o_data_a = 16'b0000000000000000;
            14'h1470: o_data_a = 16'b1111110010101000;
            14'h1471: o_data_a = 16'b1111110000010000;
            14'h1472: o_data_a = 16'b0000000000000011;
            14'h1473: o_data_a = 16'b1111110111100000;
            14'h1474: o_data_a = 16'b1110110111100000;
            14'h1475: o_data_a = 16'b1110001100001000;
            14'h1476: o_data_a = 16'b0000000000000011;
            14'h1477: o_data_a = 16'b1111110111100000;
            14'h1478: o_data_a = 16'b1110110111100000;
            14'h1479: o_data_a = 16'b1111110000010000;
            14'h147a: o_data_a = 16'b0000000000000000;
            14'h147b: o_data_a = 16'b1111110111101000;
            14'h147c: o_data_a = 16'b1110110010100000;
            14'h147d: o_data_a = 16'b1110001100001000;
            14'h147e: o_data_a = 16'b0000000000000000;
            14'h147f: o_data_a = 16'b1111110111001000;
            14'h1480: o_data_a = 16'b1111110010100000;
            14'h1481: o_data_a = 16'b1110101010001000;
            14'h1482: o_data_a = 16'b0001010010000110;
            14'h1483: o_data_a = 16'b1110110000010000;
            14'h1484: o_data_a = 16'b0000000000010110;
            14'h1485: o_data_a = 16'b1110101010000111;
            14'h1486: o_data_a = 16'b0000000000000011;
            14'h1487: o_data_a = 16'b1111110111100000;
            14'h1488: o_data_a = 16'b1110110111100000;
            14'h1489: o_data_a = 16'b1111110000010000;
            14'h148a: o_data_a = 16'b0000000000000000;
            14'h148b: o_data_a = 16'b1111110111101000;
            14'h148c: o_data_a = 16'b1110110010100000;
            14'h148d: o_data_a = 16'b1110001100001000;
            14'h148e: o_data_a = 16'b0000000000000011;
            14'h148f: o_data_a = 16'b1111110000010000;
            14'h1490: o_data_a = 16'b0000000000000101;
            14'h1491: o_data_a = 16'b1110000010100000;
            14'h1492: o_data_a = 16'b1111110000010000;
            14'h1493: o_data_a = 16'b0000000000000000;
            14'h1494: o_data_a = 16'b1111110111101000;
            14'h1495: o_data_a = 16'b1110110010100000;
            14'h1496: o_data_a = 16'b1110001100001000;
            14'h1497: o_data_a = 16'b0001010010011011;
            14'h1498: o_data_a = 16'b1110110000010000;
            14'h1499: o_data_a = 16'b0000000000000110;
            14'h149a: o_data_a = 16'b1110101010000111;
            14'h149b: o_data_a = 16'b0000000000000000;
            14'h149c: o_data_a = 16'b1111110010100000;
            14'h149d: o_data_a = 16'b1111110001001000;
            14'h149e: o_data_a = 16'b0000000000000000;
            14'h149f: o_data_a = 16'b1111110010101000;
            14'h14a0: o_data_a = 16'b1111110000010000;
            14'h14a1: o_data_a = 16'b1110110010100000;
            14'h14a2: o_data_a = 16'b1111000000001000;
            14'h14a3: o_data_a = 16'b0000000000000000;
            14'h14a4: o_data_a = 16'b1111110010101000;
            14'h14a5: o_data_a = 16'b1111110000010000;
            14'h14a6: o_data_a = 16'b0001010010101010;
            14'h14a7: o_data_a = 16'b1110001100000101;
            14'h14a8: o_data_a = 16'b0001011010101010;
            14'h14a9: o_data_a = 16'b1110101010000111;
            14'h14aa: o_data_a = 16'b0000000000000011;
            14'h14ab: o_data_a = 16'b1111110111100000;
            14'h14ac: o_data_a = 16'b1110110111100000;
            14'h14ad: o_data_a = 16'b1111110000010000;
            14'h14ae: o_data_a = 16'b0000000000000000;
            14'h14af: o_data_a = 16'b1111110111101000;
            14'h14b0: o_data_a = 16'b1110110010100000;
            14'h14b1: o_data_a = 16'b1110001100001000;
            14'h14b2: o_data_a = 16'b0000000000000000;
            14'h14b3: o_data_a = 16'b1111110010101000;
            14'h14b4: o_data_a = 16'b1111110000010000;
            14'h14b5: o_data_a = 16'b0000000000000011;
            14'h14b6: o_data_a = 16'b1111110111100000;
            14'h14b7: o_data_a = 16'b1110110111100000;
            14'h14b8: o_data_a = 16'b1110110111100000;
            14'h14b9: o_data_a = 16'b1110110111100000;
            14'h14ba: o_data_a = 16'b1110110111100000;
            14'h14bb: o_data_a = 16'b1110001100001000;
            14'h14bc: o_data_a = 16'b0000000000000000;
            14'h14bd: o_data_a = 16'b1111110111001000;
            14'h14be: o_data_a = 16'b1111110010100000;
            14'h14bf: o_data_a = 16'b1110101010001000;
            14'h14c0: o_data_a = 16'b0000000000000000;
            14'h14c1: o_data_a = 16'b1111110010101000;
            14'h14c2: o_data_a = 16'b1111110000010000;
            14'h14c3: o_data_a = 16'b0000000000000001;
            14'h14c4: o_data_a = 16'b1111110000100000;
            14'h14c5: o_data_a = 16'b1110001100001000;
            14'h14c6: o_data_a = 16'b0000000000000011;
            14'h14c7: o_data_a = 16'b1111110000100000;
            14'h14c8: o_data_a = 16'b1111110000010000;
            14'h14c9: o_data_a = 16'b0000000000000000;
            14'h14ca: o_data_a = 16'b1111110111101000;
            14'h14cb: o_data_a = 16'b1110110010100000;
            14'h14cc: o_data_a = 16'b1110001100001000;
            14'h14cd: o_data_a = 16'b0000000000000001;
            14'h14ce: o_data_a = 16'b1110110000010000;
            14'h14cf: o_data_a = 16'b0000000000001101;
            14'h14d0: o_data_a = 16'b1110001100001000;
            14'h14d1: o_data_a = 16'b0000110000000110;
            14'h14d2: o_data_a = 16'b1110110000010000;
            14'h14d3: o_data_a = 16'b0000000000001110;
            14'h14d4: o_data_a = 16'b1110001100001000;
            14'h14d5: o_data_a = 16'b0001010011011001;
            14'h14d6: o_data_a = 16'b1110110000010000;
            14'h14d7: o_data_a = 16'b0000000001011111;
            14'h14d8: o_data_a = 16'b1110101010000111;
            14'h14d9: o_data_a = 16'b0000000000000000;
            14'h14da: o_data_a = 16'b1111110010101000;
            14'h14db: o_data_a = 16'b1111110000010000;
            14'h14dc: o_data_a = 16'b0000000000000001;
            14'h14dd: o_data_a = 16'b1111110111100000;
            14'h14de: o_data_a = 16'b1110001100001000;
            14'h14df: o_data_a = 16'b0000000000000011;
            14'h14e0: o_data_a = 16'b1111110000100000;
            14'h14e1: o_data_a = 16'b1111110000010000;
            14'h14e2: o_data_a = 16'b0000000000000000;
            14'h14e3: o_data_a = 16'b1111110111101000;
            14'h14e4: o_data_a = 16'b1110110010100000;
            14'h14e5: o_data_a = 16'b1110001100001000;
            14'h14e6: o_data_a = 16'b0000000000000001;
            14'h14e7: o_data_a = 16'b1110110000010000;
            14'h14e8: o_data_a = 16'b0000000000001101;
            14'h14e9: o_data_a = 16'b1110001100001000;
            14'h14ea: o_data_a = 16'b0000110000011011;
            14'h14eb: o_data_a = 16'b1110110000010000;
            14'h14ec: o_data_a = 16'b0000000000001110;
            14'h14ed: o_data_a = 16'b1110001100001000;
            14'h14ee: o_data_a = 16'b0001010011110010;
            14'h14ef: o_data_a = 16'b1110110000010000;
            14'h14f0: o_data_a = 16'b0000000001011111;
            14'h14f1: o_data_a = 16'b1110101010000111;
            14'h14f2: o_data_a = 16'b0000000000000000;
            14'h14f3: o_data_a = 16'b1111110010101000;
            14'h14f4: o_data_a = 16'b1111110000010000;
            14'h14f5: o_data_a = 16'b0000000000000001;
            14'h14f6: o_data_a = 16'b1111110111100000;
            14'h14f7: o_data_a = 16'b1110110111100000;
            14'h14f8: o_data_a = 16'b1110001100001000;
            14'h14f9: o_data_a = 16'b0000000000000011;
            14'h14fa: o_data_a = 16'b1111110111100000;
            14'h14fb: o_data_a = 16'b1111110000010000;
            14'h14fc: o_data_a = 16'b0000000000000000;
            14'h14fd: o_data_a = 16'b1111110111101000;
            14'h14fe: o_data_a = 16'b1110110010100000;
            14'h14ff: o_data_a = 16'b1110001100001000;
            14'h1500: o_data_a = 16'b0000000000000001;
            14'h1501: o_data_a = 16'b1110110000010000;
            14'h1502: o_data_a = 16'b0000000000001101;
            14'h1503: o_data_a = 16'b1110001100001000;
            14'h1504: o_data_a = 16'b0000001001010111;
            14'h1505: o_data_a = 16'b1110110000010000;
            14'h1506: o_data_a = 16'b0000000000001110;
            14'h1507: o_data_a = 16'b1110001100001000;
            14'h1508: o_data_a = 16'b0001010100001100;
            14'h1509: o_data_a = 16'b1110110000010000;
            14'h150a: o_data_a = 16'b0000000001011111;
            14'h150b: o_data_a = 16'b1110101010000111;
            14'h150c: o_data_a = 16'b0000000000000000;
            14'h150d: o_data_a = 16'b1111110010101000;
            14'h150e: o_data_a = 16'b1111110000010000;
            14'h150f: o_data_a = 16'b0000000000000001;
            14'h1510: o_data_a = 16'b1111110111100000;
            14'h1511: o_data_a = 16'b1110110111100000;
            14'h1512: o_data_a = 16'b1110110111100000;
            14'h1513: o_data_a = 16'b1110001100001000;
            14'h1514: o_data_a = 16'b0000000000000011;
            14'h1515: o_data_a = 16'b1111110111100000;
            14'h1516: o_data_a = 16'b1111110000010000;
            14'h1517: o_data_a = 16'b0000000000000000;
            14'h1518: o_data_a = 16'b1111110111101000;
            14'h1519: o_data_a = 16'b1110110010100000;
            14'h151a: o_data_a = 16'b1110001100001000;
            14'h151b: o_data_a = 16'b0000000000000001;
            14'h151c: o_data_a = 16'b1110110000010000;
            14'h151d: o_data_a = 16'b0000000000001101;
            14'h151e: o_data_a = 16'b1110001100001000;
            14'h151f: o_data_a = 16'b0000001001101100;
            14'h1520: o_data_a = 16'b1110110000010000;
            14'h1521: o_data_a = 16'b0000000000001110;
            14'h1522: o_data_a = 16'b1110001100001000;
            14'h1523: o_data_a = 16'b0001010100100111;
            14'h1524: o_data_a = 16'b1110110000010000;
            14'h1525: o_data_a = 16'b0000000001011111;
            14'h1526: o_data_a = 16'b1110101010000111;
            14'h1527: o_data_a = 16'b0000000000000000;
            14'h1528: o_data_a = 16'b1111110010101000;
            14'h1529: o_data_a = 16'b1111110000010000;
            14'h152a: o_data_a = 16'b0000000000000001;
            14'h152b: o_data_a = 16'b1111110111100000;
            14'h152c: o_data_a = 16'b1110110111100000;
            14'h152d: o_data_a = 16'b1110110111100000;
            14'h152e: o_data_a = 16'b1110110111100000;
            14'h152f: o_data_a = 16'b1110001100001000;
            14'h1530: o_data_a = 16'b0000000000000011;
            14'h1531: o_data_a = 16'b1111110111100000;
            14'h1532: o_data_a = 16'b1110110111100000;
            14'h1533: o_data_a = 16'b1111110000010000;
            14'h1534: o_data_a = 16'b0000000000000000;
            14'h1535: o_data_a = 16'b1111110111101000;
            14'h1536: o_data_a = 16'b1110110010100000;
            14'h1537: o_data_a = 16'b1110001100001000;
            14'h1538: o_data_a = 16'b0000000000000100;
            14'h1539: o_data_a = 16'b1110110000010000;
            14'h153a: o_data_a = 16'b0000000000000000;
            14'h153b: o_data_a = 16'b1111110111101000;
            14'h153c: o_data_a = 16'b1110110010100000;
            14'h153d: o_data_a = 16'b1110001100001000;
            14'h153e: o_data_a = 16'b0001010101000010;
            14'h153f: o_data_a = 16'b1110110000010000;
            14'h1540: o_data_a = 16'b0000000000000110;
            14'h1541: o_data_a = 16'b1110101010000111;
            14'h1542: o_data_a = 16'b0000000000000000;
            14'h1543: o_data_a = 16'b1111110010101000;
            14'h1544: o_data_a = 16'b1111110000010000;
            14'h1545: o_data_a = 16'b0001010101001001;
            14'h1546: o_data_a = 16'b1110001100000101;
            14'h1547: o_data_a = 16'b0001011010001011;
            14'h1548: o_data_a = 16'b1110101010000111;
            14'h1549: o_data_a = 16'b0000000000000001;
            14'h154a: o_data_a = 16'b1111110111100000;
            14'h154b: o_data_a = 16'b1111110000010000;
            14'h154c: o_data_a = 16'b0000000000000000;
            14'h154d: o_data_a = 16'b1111110111101000;
            14'h154e: o_data_a = 16'b1110110010100000;
            14'h154f: o_data_a = 16'b1110001100001000;
            14'h1550: o_data_a = 16'b0000000000000001;
            14'h1551: o_data_a = 16'b1111110000010000;
            14'h1552: o_data_a = 16'b0000000000000100;
            14'h1553: o_data_a = 16'b1110000010100000;
            14'h1554: o_data_a = 16'b1111110000010000;
            14'h1555: o_data_a = 16'b0000000000000000;
            14'h1556: o_data_a = 16'b1111110111101000;
            14'h1557: o_data_a = 16'b1110110010100000;
            14'h1558: o_data_a = 16'b1110001100001000;
            14'h1559: o_data_a = 16'b0001010101011101;
            14'h155a: o_data_a = 16'b1110110000010000;
            14'h155b: o_data_a = 16'b0000000000010110;
            14'h155c: o_data_a = 16'b1110101010000111;
            14'h155d: o_data_a = 16'b0000000000000001;
            14'h155e: o_data_a = 16'b1111110111100000;
            14'h155f: o_data_a = 16'b1110110111100000;
            14'h1560: o_data_a = 16'b1111110000010000;
            14'h1561: o_data_a = 16'b0000000000000000;
            14'h1562: o_data_a = 16'b1111110111101000;
            14'h1563: o_data_a = 16'b1110110010100000;
            14'h1564: o_data_a = 16'b1110001100001000;
            14'h1565: o_data_a = 16'b0000000000000001;
            14'h1566: o_data_a = 16'b1111110000010000;
            14'h1567: o_data_a = 16'b0000000000000011;
            14'h1568: o_data_a = 16'b1110000010100000;
            14'h1569: o_data_a = 16'b1111110000010000;
            14'h156a: o_data_a = 16'b0000000000000000;
            14'h156b: o_data_a = 16'b1111110111101000;
            14'h156c: o_data_a = 16'b1110110010100000;
            14'h156d: o_data_a = 16'b1110001100001000;
            14'h156e: o_data_a = 16'b0001010101110010;
            14'h156f: o_data_a = 16'b1110110000010000;
            14'h1570: o_data_a = 16'b0000000000100110;
            14'h1571: o_data_a = 16'b1110101010000111;
            14'h1572: o_data_a = 16'b0000000000000000;
            14'h1573: o_data_a = 16'b1111110010101000;
            14'h1574: o_data_a = 16'b1111110000010000;
            14'h1575: o_data_a = 16'b1110110010100000;
            14'h1576: o_data_a = 16'b1111010101001000;
            14'h1577: o_data_a = 16'b0000000000000000;
            14'h1578: o_data_a = 16'b1111110010101000;
            14'h1579: o_data_a = 16'b1111110000010000;
            14'h157a: o_data_a = 16'b0000000000000011;
            14'h157b: o_data_a = 16'b1111110111100000;
            14'h157c: o_data_a = 16'b1110110111100000;
            14'h157d: o_data_a = 16'b1110110111100000;
            14'h157e: o_data_a = 16'b1110001100001000;
            14'h157f: o_data_a = 16'b0000000000000011;
            14'h1580: o_data_a = 16'b1111110000010000;
            14'h1581: o_data_a = 16'b0000000000000011;
            14'h1582: o_data_a = 16'b1110000010100000;
            14'h1583: o_data_a = 16'b1111110000010000;
            14'h1584: o_data_a = 16'b0000000000000000;
            14'h1585: o_data_a = 16'b1111110111101000;
            14'h1586: o_data_a = 16'b1110110010100000;
            14'h1587: o_data_a = 16'b1110001100001000;
            14'h1588: o_data_a = 16'b0000000000000000;
            14'h1589: o_data_a = 16'b1111110010100000;
            14'h158a: o_data_a = 16'b1111110001001000;
            14'h158b: o_data_a = 16'b0000000000000000;
            14'h158c: o_data_a = 16'b1111110010101000;
            14'h158d: o_data_a = 16'b1111110000010000;
            14'h158e: o_data_a = 16'b0001010110010010;
            14'h158f: o_data_a = 16'b1110001100000101;
            14'h1590: o_data_a = 16'b0001011010001011;
            14'h1591: o_data_a = 16'b1110101010000111;
            14'h1592: o_data_a = 16'b0000000000000001;
            14'h1593: o_data_a = 16'b1111110000010000;
            14'h1594: o_data_a = 16'b0000000000000100;
            14'h1595: o_data_a = 16'b1110000010100000;
            14'h1596: o_data_a = 16'b1111110000010000;
            14'h1597: o_data_a = 16'b0000000000000000;
            14'h1598: o_data_a = 16'b1111110111101000;
            14'h1599: o_data_a = 16'b1110110010100000;
            14'h159a: o_data_a = 16'b1110001100001000;
            14'h159b: o_data_a = 16'b0000000000000001;
            14'h159c: o_data_a = 16'b1111110111100000;
            14'h159d: o_data_a = 16'b1111110000010000;
            14'h159e: o_data_a = 16'b0000000000000000;
            14'h159f: o_data_a = 16'b1111110111101000;
            14'h15a0: o_data_a = 16'b1110110010100000;
            14'h15a1: o_data_a = 16'b1110001100001000;
            14'h15a2: o_data_a = 16'b0000000000001010;
            14'h15a3: o_data_a = 16'b1110110000010000;
            14'h15a4: o_data_a = 16'b0000000000000000;
            14'h15a5: o_data_a = 16'b1111110111101000;
            14'h15a6: o_data_a = 16'b1110110010100000;
            14'h15a7: o_data_a = 16'b1110001100001000;
            14'h15a8: o_data_a = 16'b0000000000000000;
            14'h15a9: o_data_a = 16'b1111110010101000;
            14'h15aa: o_data_a = 16'b1111110000010000;
            14'h15ab: o_data_a = 16'b1110110010100000;
            14'h15ac: o_data_a = 16'b1111000010001000;
            14'h15ad: o_data_a = 16'b0001010110110001;
            14'h15ae: o_data_a = 16'b1110110000010000;
            14'h15af: o_data_a = 16'b0000000000100110;
            14'h15b0: o_data_a = 16'b1110101010000111;
            14'h15b1: o_data_a = 16'b0000000000000000;
            14'h15b2: o_data_a = 16'b1111110010101000;
            14'h15b3: o_data_a = 16'b1111110000010000;
            14'h15b4: o_data_a = 16'b0001010110111000;
            14'h15b5: o_data_a = 16'b1110001100000101;
            14'h15b6: o_data_a = 16'b0001010111001000;
            14'h15b7: o_data_a = 16'b1110101010000111;
            14'h15b8: o_data_a = 16'b0000000000000000;
            14'h15b9: o_data_a = 16'b1111110111001000;
            14'h15ba: o_data_a = 16'b1111110010100000;
            14'h15bb: o_data_a = 16'b1110111111001000;
            14'h15bc: o_data_a = 16'b0000000000000000;
            14'h15bd: o_data_a = 16'b1111110010100000;
            14'h15be: o_data_a = 16'b1111110001010000;
            14'h15bf: o_data_a = 16'b1110011111001000;
            14'h15c0: o_data_a = 16'b0000000000000000;
            14'h15c1: o_data_a = 16'b1111110010101000;
            14'h15c2: o_data_a = 16'b1111110000010000;
            14'h15c3: o_data_a = 16'b0000000000000001;
            14'h15c4: o_data_a = 16'b1111110000100000;
            14'h15c5: o_data_a = 16'b1110001100001000;
            14'h15c6: o_data_a = 16'b0001010111111001;
            14'h15c7: o_data_a = 16'b1110101010000111;
            14'h15c8: o_data_a = 16'b0000000000000001;
            14'h15c9: o_data_a = 16'b1111110000010000;
            14'h15ca: o_data_a = 16'b0000000000000011;
            14'h15cb: o_data_a = 16'b1110000010100000;
            14'h15cc: o_data_a = 16'b1111110000010000;
            14'h15cd: o_data_a = 16'b0000000000000000;
            14'h15ce: o_data_a = 16'b1111110111101000;
            14'h15cf: o_data_a = 16'b1110110010100000;
            14'h15d0: o_data_a = 16'b1110001100001000;
            14'h15d1: o_data_a = 16'b0000000000000001;
            14'h15d2: o_data_a = 16'b1111110111100000;
            14'h15d3: o_data_a = 16'b1110110111100000;
            14'h15d4: o_data_a = 16'b1111110000010000;
            14'h15d5: o_data_a = 16'b0000000000000000;
            14'h15d6: o_data_a = 16'b1111110111101000;
            14'h15d7: o_data_a = 16'b1110110010100000;
            14'h15d8: o_data_a = 16'b1110001100001000;
            14'h15d9: o_data_a = 16'b0000000000001010;
            14'h15da: o_data_a = 16'b1110110000010000;
            14'h15db: o_data_a = 16'b0000000000000000;
            14'h15dc: o_data_a = 16'b1111110111101000;
            14'h15dd: o_data_a = 16'b1110110010100000;
            14'h15de: o_data_a = 16'b1110001100001000;
            14'h15df: o_data_a = 16'b0000000000000000;
            14'h15e0: o_data_a = 16'b1111110010101000;
            14'h15e1: o_data_a = 16'b1111110000010000;
            14'h15e2: o_data_a = 16'b1110110010100000;
            14'h15e3: o_data_a = 16'b1111000111001000;
            14'h15e4: o_data_a = 16'b0001010111101000;
            14'h15e5: o_data_a = 16'b1110110000010000;
            14'h15e6: o_data_a = 16'b0000000000010110;
            14'h15e7: o_data_a = 16'b1110101010000111;
            14'h15e8: o_data_a = 16'b0000000000000000;
            14'h15e9: o_data_a = 16'b1111110010101000;
            14'h15ea: o_data_a = 16'b1111110000010000;
            14'h15eb: o_data_a = 16'b0001010111101111;
            14'h15ec: o_data_a = 16'b1110001100000101;
            14'h15ed: o_data_a = 16'b0001010111111001;
            14'h15ee: o_data_a = 16'b1110101010000111;
            14'h15ef: o_data_a = 16'b0000000000000000;
            14'h15f0: o_data_a = 16'b1111110111001000;
            14'h15f1: o_data_a = 16'b1111110010100000;
            14'h15f2: o_data_a = 16'b1110111111001000;
            14'h15f3: o_data_a = 16'b0000000000000000;
            14'h15f4: o_data_a = 16'b1111110010101000;
            14'h15f5: o_data_a = 16'b1111110000010000;
            14'h15f6: o_data_a = 16'b0000000000000001;
            14'h15f7: o_data_a = 16'b1111110000100000;
            14'h15f8: o_data_a = 16'b1110001100001000;
            14'h15f9: o_data_a = 16'b0000000000000011;
            14'h15fa: o_data_a = 16'b1111110000010000;
            14'h15fb: o_data_a = 16'b0000000000000110;
            14'h15fc: o_data_a = 16'b1110000010100000;
            14'h15fd: o_data_a = 16'b1111110000010000;
            14'h15fe: o_data_a = 16'b0000000000000000;
            14'h15ff: o_data_a = 16'b1111110111101000;
            14'h1600: o_data_a = 16'b1110110010100000;
            14'h1601: o_data_a = 16'b1110001100001000;
            14'h1602: o_data_a = 16'b0000000000000010;
            14'h1603: o_data_a = 16'b1110110000010000;
            14'h1604: o_data_a = 16'b0000000000000000;
            14'h1605: o_data_a = 16'b1111110111101000;
            14'h1606: o_data_a = 16'b1110110010100000;
            14'h1607: o_data_a = 16'b1110001100001000;
            14'h1608: o_data_a = 16'b0000000000000000;
            14'h1609: o_data_a = 16'b1111110010101000;
            14'h160a: o_data_a = 16'b1111110000010000;
            14'h160b: o_data_a = 16'b1110110010100000;
            14'h160c: o_data_a = 16'b1111000111001000;
            14'h160d: o_data_a = 16'b0000000000000000;
            14'h160e: o_data_a = 16'b1111110010101000;
            14'h160f: o_data_a = 16'b1111110000010000;
            14'h1610: o_data_a = 16'b0000000000000011;
            14'h1611: o_data_a = 16'b1111110111100000;
            14'h1612: o_data_a = 16'b1110110111100000;
            14'h1613: o_data_a = 16'b1110110111100000;
            14'h1614: o_data_a = 16'b1110110111100000;
            14'h1615: o_data_a = 16'b1110110111100000;
            14'h1616: o_data_a = 16'b1110110111100000;
            14'h1617: o_data_a = 16'b1110001100001000;
            14'h1618: o_data_a = 16'b0000000000000011;
            14'h1619: o_data_a = 16'b1111110000100000;
            14'h161a: o_data_a = 16'b1111110000010000;
            14'h161b: o_data_a = 16'b0000000000000000;
            14'h161c: o_data_a = 16'b1111110111101000;
            14'h161d: o_data_a = 16'b1110110010100000;
            14'h161e: o_data_a = 16'b1110001100001000;
            14'h161f: o_data_a = 16'b0000000000000011;
            14'h1620: o_data_a = 16'b1111110000010000;
            14'h1621: o_data_a = 16'b0000000000000110;
            14'h1622: o_data_a = 16'b1110000010100000;
            14'h1623: o_data_a = 16'b1111110000010000;
            14'h1624: o_data_a = 16'b0000000000000000;
            14'h1625: o_data_a = 16'b1111110111101000;
            14'h1626: o_data_a = 16'b1110110010100000;
            14'h1627: o_data_a = 16'b1110001100001000;
            14'h1628: o_data_a = 16'b0000000000000010;
            14'h1629: o_data_a = 16'b1110110000010000;
            14'h162a: o_data_a = 16'b0000000000001101;
            14'h162b: o_data_a = 16'b1110001100001000;
            14'h162c: o_data_a = 16'b0000110000111101;
            14'h162d: o_data_a = 16'b1110110000010000;
            14'h162e: o_data_a = 16'b0000000000001110;
            14'h162f: o_data_a = 16'b1110001100001000;
            14'h1630: o_data_a = 16'b0001011000110100;
            14'h1631: o_data_a = 16'b1110110000010000;
            14'h1632: o_data_a = 16'b0000000001011111;
            14'h1633: o_data_a = 16'b1110101010000111;
            14'h1634: o_data_a = 16'b0000000000000000;
            14'h1635: o_data_a = 16'b1111110010101000;
            14'h1636: o_data_a = 16'b1111110000010000;
            14'h1637: o_data_a = 16'b0000000000000101;
            14'h1638: o_data_a = 16'b1110001100001000;
            14'h1639: o_data_a = 16'b0000000000000011;
            14'h163a: o_data_a = 16'b1111110000010000;
            14'h163b: o_data_a = 16'b0000000000000100;
            14'h163c: o_data_a = 16'b1110000010100000;
            14'h163d: o_data_a = 16'b1111110000010000;
            14'h163e: o_data_a = 16'b0000000000000000;
            14'h163f: o_data_a = 16'b1111110111101000;
            14'h1640: o_data_a = 16'b1110110010100000;
            14'h1641: o_data_a = 16'b1110001100001000;
            14'h1642: o_data_a = 16'b0000000000000000;
            14'h1643: o_data_a = 16'b1111110111001000;
            14'h1644: o_data_a = 16'b1111110010100000;
            14'h1645: o_data_a = 16'b1110111111001000;
            14'h1646: o_data_a = 16'b0000000000000000;
            14'h1647: o_data_a = 16'b1111110010101000;
            14'h1648: o_data_a = 16'b1111110000010000;
            14'h1649: o_data_a = 16'b1110110010100000;
            14'h164a: o_data_a = 16'b1111000010001000;
            14'h164b: o_data_a = 16'b0000000000000000;
            14'h164c: o_data_a = 16'b1111110010101000;
            14'h164d: o_data_a = 16'b1111110000010000;
            14'h164e: o_data_a = 16'b0000000000000011;
            14'h164f: o_data_a = 16'b1111110111100000;
            14'h1650: o_data_a = 16'b1110110111100000;
            14'h1651: o_data_a = 16'b1110110111100000;
            14'h1652: o_data_a = 16'b1110110111100000;
            14'h1653: o_data_a = 16'b1110001100001000;
            14'h1654: o_data_a = 16'b0000000000010110;
            14'h1655: o_data_a = 16'b1110110000010000;
            14'h1656: o_data_a = 16'b0000000000000000;
            14'h1657: o_data_a = 16'b1111110111101000;
            14'h1658: o_data_a = 16'b1110110010100000;
            14'h1659: o_data_a = 16'b1110001100001000;
            14'h165a: o_data_a = 16'b0000000000000111;
            14'h165b: o_data_a = 16'b1110110000010000;
            14'h165c: o_data_a = 16'b0000000000000000;
            14'h165d: o_data_a = 16'b1111110111101000;
            14'h165e: o_data_a = 16'b1110110010100000;
            14'h165f: o_data_a = 16'b1110001100001000;
            14'h1660: o_data_a = 16'b0000000000000010;
            14'h1661: o_data_a = 16'b1110110000010000;
            14'h1662: o_data_a = 16'b0000000000001101;
            14'h1663: o_data_a = 16'b1110001100001000;
            14'h1664: o_data_a = 16'b0100101110010110;
            14'h1665: o_data_a = 16'b1110110000010000;
            14'h1666: o_data_a = 16'b0000000000001110;
            14'h1667: o_data_a = 16'b1110001100001000;
            14'h1668: o_data_a = 16'b0001011001101100;
            14'h1669: o_data_a = 16'b1110110000010000;
            14'h166a: o_data_a = 16'b0000000001011111;
            14'h166b: o_data_a = 16'b1110101010000111;
            14'h166c: o_data_a = 16'b0000000000000000;
            14'h166d: o_data_a = 16'b1111110010101000;
            14'h166e: o_data_a = 16'b1111110000010000;
            14'h166f: o_data_a = 16'b0000000000000101;
            14'h1670: o_data_a = 16'b1110001100001000;
            14'h1671: o_data_a = 16'b0000000000000011;
            14'h1672: o_data_a = 16'b1111110000010000;
            14'h1673: o_data_a = 16'b0000000000000100;
            14'h1674: o_data_a = 16'b1110000010100000;
            14'h1675: o_data_a = 16'b1111110000010000;
            14'h1676: o_data_a = 16'b0000000000000000;
            14'h1677: o_data_a = 16'b1111110111101000;
            14'h1678: o_data_a = 16'b1110110010100000;
            14'h1679: o_data_a = 16'b1110001100001000;
            14'h167a: o_data_a = 16'b0000000000000001;
            14'h167b: o_data_a = 16'b1110110000010000;
            14'h167c: o_data_a = 16'b0000000000001101;
            14'h167d: o_data_a = 16'b1110001100001000;
            14'h167e: o_data_a = 16'b0100111000001101;
            14'h167f: o_data_a = 16'b1110110000010000;
            14'h1680: o_data_a = 16'b0000000000001110;
            14'h1681: o_data_a = 16'b1110001100001000;
            14'h1682: o_data_a = 16'b0001011010000110;
            14'h1683: o_data_a = 16'b1110110000010000;
            14'h1684: o_data_a = 16'b0000000001011111;
            14'h1685: o_data_a = 16'b1110101010000111;
            14'h1686: o_data_a = 16'b0000000000000000;
            14'h1687: o_data_a = 16'b1111110010101000;
            14'h1688: o_data_a = 16'b1111110000010000;
            14'h1689: o_data_a = 16'b0000000000000101;
            14'h168a: o_data_a = 16'b1110001100001000;
            14'h168b: o_data_a = 16'b0000000000000011;
            14'h168c: o_data_a = 16'b1111110111100000;
            14'h168d: o_data_a = 16'b1111110000010000;
            14'h168e: o_data_a = 16'b0000000000000000;
            14'h168f: o_data_a = 16'b1111110111101000;
            14'h1690: o_data_a = 16'b1110110010100000;
            14'h1691: o_data_a = 16'b1110001100001000;
            14'h1692: o_data_a = 16'b0000000000000001;
            14'h1693: o_data_a = 16'b1111110000100000;
            14'h1694: o_data_a = 16'b1111110000010000;
            14'h1695: o_data_a = 16'b0000000000000000;
            14'h1696: o_data_a = 16'b1111110111101000;
            14'h1697: o_data_a = 16'b1110110010100000;
            14'h1698: o_data_a = 16'b1110001100001000;
            14'h1699: o_data_a = 16'b0000000000000010;
            14'h169a: o_data_a = 16'b1110110000010000;
            14'h169b: o_data_a = 16'b0000000000001101;
            14'h169c: o_data_a = 16'b1110001100001000;
            14'h169d: o_data_a = 16'b0000011100101011;
            14'h169e: o_data_a = 16'b1110110000010000;
            14'h169f: o_data_a = 16'b0000000000001110;
            14'h16a0: o_data_a = 16'b1110001100001000;
            14'h16a1: o_data_a = 16'b0001011010100101;
            14'h16a2: o_data_a = 16'b1110110000010000;
            14'h16a3: o_data_a = 16'b0000000001011111;
            14'h16a4: o_data_a = 16'b1110101010000111;
            14'h16a5: o_data_a = 16'b0000000000000000;
            14'h16a6: o_data_a = 16'b1111110010101000;
            14'h16a7: o_data_a = 16'b1111110000010000;
            14'h16a8: o_data_a = 16'b0000000000000101;
            14'h16a9: o_data_a = 16'b1110001100001000;
            14'h16aa: o_data_a = 16'b0000000000000000;
            14'h16ab: o_data_a = 16'b1111110111001000;
            14'h16ac: o_data_a = 16'b1111110010100000;
            14'h16ad: o_data_a = 16'b1110101010001000;
            14'h16ae: o_data_a = 16'b0000000000110110;
            14'h16af: o_data_a = 16'b1110101010000111;
            14'h16b0: o_data_a = 16'b0000000000000010;
            14'h16b1: o_data_a = 16'b1111110000100000;
            14'h16b2: o_data_a = 16'b1111110000010000;
            14'h16b3: o_data_a = 16'b0000000000000000;
            14'h16b4: o_data_a = 16'b1111110111101000;
            14'h16b5: o_data_a = 16'b1110110010100000;
            14'h16b6: o_data_a = 16'b1110001100001000;
            14'h16b7: o_data_a = 16'b0000000000000000;
            14'h16b8: o_data_a = 16'b1111110111001000;
            14'h16b9: o_data_a = 16'b1111110010100000;
            14'h16ba: o_data_a = 16'b1110101010001000;
            14'h16bb: o_data_a = 16'b0001011010111111;
            14'h16bc: o_data_a = 16'b1110110000010000;
            14'h16bd: o_data_a = 16'b0000000000010110;
            14'h16be: o_data_a = 16'b1110101010000111;
            14'h16bf: o_data_a = 16'b0000000000000000;
            14'h16c0: o_data_a = 16'b1111110010100000;
            14'h16c1: o_data_a = 16'b1111110001001000;
            14'h16c2: o_data_a = 16'b0000000000000000;
            14'h16c3: o_data_a = 16'b1111110010101000;
            14'h16c4: o_data_a = 16'b1111110000010000;
            14'h16c5: o_data_a = 16'b0001011011001001;
            14'h16c6: o_data_a = 16'b1110001100000101;
            14'h16c7: o_data_a = 16'b0001011011100000;
            14'h16c8: o_data_a = 16'b1110101010000111;
            14'h16c9: o_data_a = 16'b0000000000000010;
            14'h16ca: o_data_a = 16'b1110110000010000;
            14'h16cb: o_data_a = 16'b0000000000000000;
            14'h16cc: o_data_a = 16'b1111110111101000;
            14'h16cd: o_data_a = 16'b1110110010100000;
            14'h16ce: o_data_a = 16'b1110001100001000;
            14'h16cf: o_data_a = 16'b0000000000000001;
            14'h16d0: o_data_a = 16'b1110110000010000;
            14'h16d1: o_data_a = 16'b0000000000001101;
            14'h16d2: o_data_a = 16'b1110001100001000;
            14'h16d3: o_data_a = 16'b0110101011011001;
            14'h16d4: o_data_a = 16'b1110110000010000;
            14'h16d5: o_data_a = 16'b0000000000001110;
            14'h16d6: o_data_a = 16'b1110001100001000;
            14'h16d7: o_data_a = 16'b0001011011011011;
            14'h16d8: o_data_a = 16'b1110110000010000;
            14'h16d9: o_data_a = 16'b0000000001011111;
            14'h16da: o_data_a = 16'b1110101010000111;
            14'h16db: o_data_a = 16'b0000000000000000;
            14'h16dc: o_data_a = 16'b1111110010101000;
            14'h16dd: o_data_a = 16'b1111110000010000;
            14'h16de: o_data_a = 16'b0000000000000101;
            14'h16df: o_data_a = 16'b1110001100001000;
            14'h16e0: o_data_a = 16'b0000000000000010;
            14'h16e1: o_data_a = 16'b1111110000100000;
            14'h16e2: o_data_a = 16'b1111110000010000;
            14'h16e3: o_data_a = 16'b0000000000000000;
            14'h16e4: o_data_a = 16'b1111110111101000;
            14'h16e5: o_data_a = 16'b1110110010100000;
            14'h16e6: o_data_a = 16'b1110001100001000;
            14'h16e7: o_data_a = 16'b0000000000000001;
            14'h16e8: o_data_a = 16'b1110110000010000;
            14'h16e9: o_data_a = 16'b0000000000001101;
            14'h16ea: o_data_a = 16'b1110001100001000;
            14'h16eb: o_data_a = 16'b0010000111000011;
            14'h16ec: o_data_a = 16'b1110110000010000;
            14'h16ed: o_data_a = 16'b0000000000001110;
            14'h16ee: o_data_a = 16'b1110001100001000;
            14'h16ef: o_data_a = 16'b0001011011110011;
            14'h16f0: o_data_a = 16'b1110110000010000;
            14'h16f1: o_data_a = 16'b0000000001011111;
            14'h16f2: o_data_a = 16'b1110101010000111;
            14'h16f3: o_data_a = 16'b0000000000110110;
            14'h16f4: o_data_a = 16'b1110101010000111;
            14'h16f5: o_data_a = 16'b0000000000000010;
            14'h16f6: o_data_a = 16'b1111110000100000;
            14'h16f7: o_data_a = 16'b1111110000010000;
            14'h16f8: o_data_a = 16'b0000000000000000;
            14'h16f9: o_data_a = 16'b1111110111101000;
            14'h16fa: o_data_a = 16'b1110110010100000;
            14'h16fb: o_data_a = 16'b1110001100001000;
            14'h16fc: o_data_a = 16'b0000000000000000;
            14'h16fd: o_data_a = 16'b1111110010101000;
            14'h16fe: o_data_a = 16'b1111110000010000;
            14'h16ff: o_data_a = 16'b0000000000000011;
            14'h1700: o_data_a = 16'b1110001100001000;
            14'h1701: o_data_a = 16'b0000000000000011;
            14'h1702: o_data_a = 16'b1111110000010000;
            14'h1703: o_data_a = 16'b0000000000000000;
            14'h1704: o_data_a = 16'b1111110111101000;
            14'h1705: o_data_a = 16'b1110110010100000;
            14'h1706: o_data_a = 16'b1110001100001000;
            14'h1707: o_data_a = 16'b0000000000000001;
            14'h1708: o_data_a = 16'b1110110000010000;
            14'h1709: o_data_a = 16'b0000000000001101;
            14'h170a: o_data_a = 16'b1110001100001000;
            14'h170b: o_data_a = 16'b0010010010001101;
            14'h170c: o_data_a = 16'b1110110000010000;
            14'h170d: o_data_a = 16'b0000000000001110;
            14'h170e: o_data_a = 16'b1110001100001000;
            14'h170f: o_data_a = 16'b0001011100010011;
            14'h1710: o_data_a = 16'b1110110000010000;
            14'h1711: o_data_a = 16'b0000000001011111;
            14'h1712: o_data_a = 16'b1110101010000111;
            14'h1713: o_data_a = 16'b0000000000000000;
            14'h1714: o_data_a = 16'b1111110010101000;
            14'h1715: o_data_a = 16'b1111110000010000;
            14'h1716: o_data_a = 16'b0000000000000101;
            14'h1717: o_data_a = 16'b1110001100001000;
            14'h1718: o_data_a = 16'b0000000000000000;
            14'h1719: o_data_a = 16'b1111110111001000;
            14'h171a: o_data_a = 16'b1111110010100000;
            14'h171b: o_data_a = 16'b1110101010001000;
            14'h171c: o_data_a = 16'b0000000000110110;
            14'h171d: o_data_a = 16'b1110101010000111;
            14'h171e: o_data_a = 16'b0000000000000000;
            14'h171f: o_data_a = 16'b1111110111001000;
            14'h1720: o_data_a = 16'b1111110010100000;
            14'h1721: o_data_a = 16'b1110101010001000;
            14'h1722: o_data_a = 16'b0000000000110110;
            14'h1723: o_data_a = 16'b1110101010000111;
            14'h1724: o_data_a = 16'b0110000000000000;
            14'h1725: o_data_a = 16'b1110110000010000;
            14'h1726: o_data_a = 16'b0000000000000000;
            14'h1727: o_data_a = 16'b1111110111101000;
            14'h1728: o_data_a = 16'b1110110010100000;
            14'h1729: o_data_a = 16'b1110001100001000;
            14'h172a: o_data_a = 16'b0000000000000001;
            14'h172b: o_data_a = 16'b1110110000010000;
            14'h172c: o_data_a = 16'b0000000000001101;
            14'h172d: o_data_a = 16'b1110001100001000;
            14'h172e: o_data_a = 16'b0010000101101110;
            14'h172f: o_data_a = 16'b1110110000010000;
            14'h1730: o_data_a = 16'b0000000000001110;
            14'h1731: o_data_a = 16'b1110001100001000;
            14'h1732: o_data_a = 16'b0001011100110110;
            14'h1733: o_data_a = 16'b1110110000010000;
            14'h1734: o_data_a = 16'b0000000001011111;
            14'h1735: o_data_a = 16'b1110101010000111;
            14'h1736: o_data_a = 16'b0000000000110110;
            14'h1737: o_data_a = 16'b1110101010000111;
            14'h1738: o_data_a = 16'b0000000000000000;
            14'h1739: o_data_a = 16'b1111110000100000;
            14'h173a: o_data_a = 16'b1110101010001000;
            14'h173b: o_data_a = 16'b1110110111110000;
            14'h173c: o_data_a = 16'b1110101010001000;
            14'h173d: o_data_a = 16'b0000000000000000;
            14'h173e: o_data_a = 16'b1110011111001000;
            14'h173f: o_data_a = 16'b0000000000000000;
            14'h1740: o_data_a = 16'b1111110111001000;
            14'h1741: o_data_a = 16'b1111110010100000;
            14'h1742: o_data_a = 16'b1110101010001000;
            14'h1743: o_data_a = 16'b0000000000000001;
            14'h1744: o_data_a = 16'b1110110000010000;
            14'h1745: o_data_a = 16'b0000000000001101;
            14'h1746: o_data_a = 16'b1110001100001000;
            14'h1747: o_data_a = 16'b0100110010011010;
            14'h1748: o_data_a = 16'b1110110000010000;
            14'h1749: o_data_a = 16'b0000000000001110;
            14'h174a: o_data_a = 16'b1110001100001000;
            14'h174b: o_data_a = 16'b0001011101001111;
            14'h174c: o_data_a = 16'b1110110000010000;
            14'h174d: o_data_a = 16'b0000000001011111;
            14'h174e: o_data_a = 16'b1110101010000111;
            14'h174f: o_data_a = 16'b0000000000000000;
            14'h1750: o_data_a = 16'b1111110010101000;
            14'h1751: o_data_a = 16'b1111110000010000;
            14'h1752: o_data_a = 16'b0000000000000101;
            14'h1753: o_data_a = 16'b1110001100001000;
            14'h1754: o_data_a = 16'b0000000000000001;
            14'h1755: o_data_a = 16'b1111110111100000;
            14'h1756: o_data_a = 16'b1111110000010000;
            14'h1757: o_data_a = 16'b0000000000000000;
            14'h1758: o_data_a = 16'b1111110111101000;
            14'h1759: o_data_a = 16'b1110110010100000;
            14'h175a: o_data_a = 16'b1110001100001000;
            14'h175b: o_data_a = 16'b0000000000000000;
            14'h175c: o_data_a = 16'b1111110111001000;
            14'h175d: o_data_a = 16'b1111110010100000;
            14'h175e: o_data_a = 16'b1110101010001000;
            14'h175f: o_data_a = 16'b0001011101100011;
            14'h1760: o_data_a = 16'b1110110000010000;
            14'h1761: o_data_a = 16'b0000000000000110;
            14'h1762: o_data_a = 16'b1110101010000111;
            14'h1763: o_data_a = 16'b0000000000000001;
            14'h1764: o_data_a = 16'b1111110000100000;
            14'h1765: o_data_a = 16'b1111110000010000;
            14'h1766: o_data_a = 16'b0000000000000000;
            14'h1767: o_data_a = 16'b1111110111101000;
            14'h1768: o_data_a = 16'b1110110010100000;
            14'h1769: o_data_a = 16'b1110001100001000;
            14'h176a: o_data_a = 16'b0000000000000000;
            14'h176b: o_data_a = 16'b1111110111001000;
            14'h176c: o_data_a = 16'b1111110010100000;
            14'h176d: o_data_a = 16'b1110101010001000;
            14'h176e: o_data_a = 16'b0001011101110010;
            14'h176f: o_data_a = 16'b1110110000010000;
            14'h1770: o_data_a = 16'b0000000000010110;
            14'h1771: o_data_a = 16'b1110101010000111;
            14'h1772: o_data_a = 16'b0000000000000000;
            14'h1773: o_data_a = 16'b1111110010101000;
            14'h1774: o_data_a = 16'b1111110000010000;
            14'h1775: o_data_a = 16'b1110110010100000;
            14'h1776: o_data_a = 16'b1111010101001000;
            14'h1777: o_data_a = 16'b0000000000000000;
            14'h1778: o_data_a = 16'b1111110010100000;
            14'h1779: o_data_a = 16'b1111110001001000;
            14'h177a: o_data_a = 16'b0000000000000000;
            14'h177b: o_data_a = 16'b1111110010101000;
            14'h177c: o_data_a = 16'b1111110000010000;
            14'h177d: o_data_a = 16'b0001011110110110;
            14'h177e: o_data_a = 16'b1110001100000101;
            14'h177f: o_data_a = 16'b0000000000000000;
            14'h1780: o_data_a = 16'b1110110000010000;
            14'h1781: o_data_a = 16'b0000000000001101;
            14'h1782: o_data_a = 16'b1110001100001000;
            14'h1783: o_data_a = 16'b0001011100100100;
            14'h1784: o_data_a = 16'b1110110000010000;
            14'h1785: o_data_a = 16'b0000000000001110;
            14'h1786: o_data_a = 16'b1110001100001000;
            14'h1787: o_data_a = 16'b0001011110001011;
            14'h1788: o_data_a = 16'b1110110000010000;
            14'h1789: o_data_a = 16'b0000000001011111;
            14'h178a: o_data_a = 16'b1110101010000111;
            14'h178b: o_data_a = 16'b0000000000000000;
            14'h178c: o_data_a = 16'b1111110010101000;
            14'h178d: o_data_a = 16'b1111110000010000;
            14'h178e: o_data_a = 16'b0000000000000001;
            14'h178f: o_data_a = 16'b1111110000100000;
            14'h1790: o_data_a = 16'b1110001100001000;
            14'h1791: o_data_a = 16'b0000000000000001;
            14'h1792: o_data_a = 16'b1111110000100000;
            14'h1793: o_data_a = 16'b1111110000010000;
            14'h1794: o_data_a = 16'b0000000000000000;
            14'h1795: o_data_a = 16'b1111110111101000;
            14'h1796: o_data_a = 16'b1110110010100000;
            14'h1797: o_data_a = 16'b1110001100001000;
            14'h1798: o_data_a = 16'b0000000000000000;
            14'h1799: o_data_a = 16'b1111110111001000;
            14'h179a: o_data_a = 16'b1111110010100000;
            14'h179b: o_data_a = 16'b1110101010001000;
            14'h179c: o_data_a = 16'b0001011110100000;
            14'h179d: o_data_a = 16'b1110110000010000;
            14'h179e: o_data_a = 16'b0000000000010110;
            14'h179f: o_data_a = 16'b1110101010000111;
            14'h17a0: o_data_a = 16'b0000000000000000;
            14'h17a1: o_data_a = 16'b1111110010101000;
            14'h17a2: o_data_a = 16'b1111110000010000;
            14'h17a3: o_data_a = 16'b0001011110100111;
            14'h17a4: o_data_a = 16'b1110001100000101;
            14'h17a5: o_data_a = 16'b0001011110110100;
            14'h17a6: o_data_a = 16'b1110101010000111;
            14'h17a7: o_data_a = 16'b0000000000000001;
            14'h17a8: o_data_a = 16'b1111110000100000;
            14'h17a9: o_data_a = 16'b1111110000010000;
            14'h17aa: o_data_a = 16'b0000000000000000;
            14'h17ab: o_data_a = 16'b1111110111101000;
            14'h17ac: o_data_a = 16'b1110110010100000;
            14'h17ad: o_data_a = 16'b1110001100001000;
            14'h17ae: o_data_a = 16'b0000000000000000;
            14'h17af: o_data_a = 16'b1111110010101000;
            14'h17b0: o_data_a = 16'b1111110000010000;
            14'h17b1: o_data_a = 16'b0000000000000001;
            14'h17b2: o_data_a = 16'b1111110111100000;
            14'h17b3: o_data_a = 16'b1110001100001000;
            14'h17b4: o_data_a = 16'b0001011101010100;
            14'h17b5: o_data_a = 16'b1110101010000111;
            14'h17b6: o_data_a = 16'b0000000000000000;
            14'h17b7: o_data_a = 16'b1110110000010000;
            14'h17b8: o_data_a = 16'b0000000000001101;
            14'h17b9: o_data_a = 16'b1110001100001000;
            14'h17ba: o_data_a = 16'b0110100110100010;
            14'h17bb: o_data_a = 16'b1110110000010000;
            14'h17bc: o_data_a = 16'b0000000000001110;
            14'h17bd: o_data_a = 16'b1110001100001000;
            14'h17be: o_data_a = 16'b0001011111000010;
            14'h17bf: o_data_a = 16'b1110110000010000;
            14'h17c0: o_data_a = 16'b0000000001011111;
            14'h17c1: o_data_a = 16'b1110101010000111;
            14'h17c2: o_data_a = 16'b0000000000000001;
            14'h17c3: o_data_a = 16'b1110110000010000;
            14'h17c4: o_data_a = 16'b0000000000001101;
            14'h17c5: o_data_a = 16'b1110001100001000;
            14'h17c6: o_data_a = 16'b0100110010011010;
            14'h17c7: o_data_a = 16'b1110110000010000;
            14'h17c8: o_data_a = 16'b0000000000001110;
            14'h17c9: o_data_a = 16'b1110001100001000;
            14'h17ca: o_data_a = 16'b0001011111001110;
            14'h17cb: o_data_a = 16'b1110110000010000;
            14'h17cc: o_data_a = 16'b0000000001011111;
            14'h17cd: o_data_a = 16'b1110101010000111;
            14'h17ce: o_data_a = 16'b0000000000000000;
            14'h17cf: o_data_a = 16'b1111110010101000;
            14'h17d0: o_data_a = 16'b1111110000010000;
            14'h17d1: o_data_a = 16'b0000000000000101;
            14'h17d2: o_data_a = 16'b1110001100001000;
            14'h17d3: o_data_a = 16'b0000000000000001;
            14'h17d4: o_data_a = 16'b1111110111100000;
            14'h17d5: o_data_a = 16'b1111110000010000;
            14'h17d6: o_data_a = 16'b0000000000000000;
            14'h17d7: o_data_a = 16'b1111110111101000;
            14'h17d8: o_data_a = 16'b1110110010100000;
            14'h17d9: o_data_a = 16'b1110001100001000;
            14'h17da: o_data_a = 16'b0000000000000001;
            14'h17db: o_data_a = 16'b1110110000010000;
            14'h17dc: o_data_a = 16'b0000000000001101;
            14'h17dd: o_data_a = 16'b1110001100001000;
            14'h17de: o_data_a = 16'b0100110010011010;
            14'h17df: o_data_a = 16'b1110110000010000;
            14'h17e0: o_data_a = 16'b0000000000001110;
            14'h17e1: o_data_a = 16'b1110001100001000;
            14'h17e2: o_data_a = 16'b0001011111100110;
            14'h17e3: o_data_a = 16'b1110110000010000;
            14'h17e4: o_data_a = 16'b0000000001011111;
            14'h17e5: o_data_a = 16'b1110101010000111;
            14'h17e6: o_data_a = 16'b0000000000000000;
            14'h17e7: o_data_a = 16'b1111110010101000;
            14'h17e8: o_data_a = 16'b1111110000010000;
            14'h17e9: o_data_a = 16'b0000000000000101;
            14'h17ea: o_data_a = 16'b1110001100001000;
            14'h17eb: o_data_a = 16'b0000000000000001;
            14'h17ec: o_data_a = 16'b1111110111100000;
            14'h17ed: o_data_a = 16'b1111110000010000;
            14'h17ee: o_data_a = 16'b0000000000000000;
            14'h17ef: o_data_a = 16'b1111110111101000;
            14'h17f0: o_data_a = 16'b1110110010100000;
            14'h17f1: o_data_a = 16'b1110001100001000;
            14'h17f2: o_data_a = 16'b0000000000110110;
            14'h17f3: o_data_a = 16'b1110101010000111;
            14'h17f4: o_data_a = 16'b0000000000000101;
            14'h17f5: o_data_a = 16'b1110110000010000;
            14'h17f6: o_data_a = 16'b1110001110010000;
            14'h17f7: o_data_a = 16'b0000000000000000;
            14'h17f8: o_data_a = 16'b1111110111101000;
            14'h17f9: o_data_a = 16'b1110110010100000;
            14'h17fa: o_data_a = 16'b1110101010001000;
            14'h17fb: o_data_a = 16'b0001011111110110;
            14'h17fc: o_data_a = 16'b1110001100000001;
            14'h17fd: o_data_a = 16'b0000000001010000;
            14'h17fe: o_data_a = 16'b1110110000010000;
            14'h17ff: o_data_a = 16'b0000000000000000;
            14'h1800: o_data_a = 16'b1111110111101000;
            14'h1801: o_data_a = 16'b1110110010100000;
            14'h1802: o_data_a = 16'b1110001100001000;
            14'h1803: o_data_a = 16'b0000000000000001;
            14'h1804: o_data_a = 16'b1110110000010000;
            14'h1805: o_data_a = 16'b0000000000001101;
            14'h1806: o_data_a = 16'b1110001100001000;
            14'h1807: o_data_a = 16'b0110001000010001;
            14'h1808: o_data_a = 16'b1110110000010000;
            14'h1809: o_data_a = 16'b0000000000001110;
            14'h180a: o_data_a = 16'b1110001100001000;
            14'h180b: o_data_a = 16'b0001100000001111;
            14'h180c: o_data_a = 16'b1110110000010000;
            14'h180d: o_data_a = 16'b0000000001011111;
            14'h180e: o_data_a = 16'b1110101010000111;
            14'h180f: o_data_a = 16'b0000000000000000;
            14'h1810: o_data_a = 16'b1111110010101000;
            14'h1811: o_data_a = 16'b1111110000010000;
            14'h1812: o_data_a = 16'b0000000000000001;
            14'h1813: o_data_a = 16'b1111110111100000;
            14'h1814: o_data_a = 16'b1110110111100000;
            14'h1815: o_data_a = 16'b1110110111100000;
            14'h1816: o_data_a = 16'b1110001100001000;
            14'h1817: o_data_a = 16'b0000000000000010;
            14'h1818: o_data_a = 16'b1111110000100000;
            14'h1819: o_data_a = 16'b1111110000010000;
            14'h181a: o_data_a = 16'b0000000000000000;
            14'h181b: o_data_a = 16'b1111110111101000;
            14'h181c: o_data_a = 16'b1110110010100000;
            14'h181d: o_data_a = 16'b1110001100001000;
            14'h181e: o_data_a = 16'b0000000000000001;
            14'h181f: o_data_a = 16'b1110110000010000;
            14'h1820: o_data_a = 16'b0000000000001101;
            14'h1821: o_data_a = 16'b1110001100001000;
            14'h1822: o_data_a = 16'b0100110110001010;
            14'h1823: o_data_a = 16'b1110110000010000;
            14'h1824: o_data_a = 16'b0000000000001110;
            14'h1825: o_data_a = 16'b1110001100001000;
            14'h1826: o_data_a = 16'b0001100000101010;
            14'h1827: o_data_a = 16'b1110110000010000;
            14'h1828: o_data_a = 16'b0000000001011111;
            14'h1829: o_data_a = 16'b1110101010000111;
            14'h182a: o_data_a = 16'b0000000000000000;
            14'h182b: o_data_a = 16'b1111110010101000;
            14'h182c: o_data_a = 16'b1111110000010000;
            14'h182d: o_data_a = 16'b0000000000000101;
            14'h182e: o_data_a = 16'b1110001100001000;
            14'h182f: o_data_a = 16'b0000000000000000;
            14'h1830: o_data_a = 16'b1110110000010000;
            14'h1831: o_data_a = 16'b0000000000001101;
            14'h1832: o_data_a = 16'b1110001100001000;
            14'h1833: o_data_a = 16'b0110100110011010;
            14'h1834: o_data_a = 16'b1110110000010000;
            14'h1835: o_data_a = 16'b0000000000001110;
            14'h1836: o_data_a = 16'b1110001100001000;
            14'h1837: o_data_a = 16'b0001100000111011;
            14'h1838: o_data_a = 16'b1110110000010000;
            14'h1839: o_data_a = 16'b0000000001011111;
            14'h183a: o_data_a = 16'b1110101010000111;
            14'h183b: o_data_a = 16'b0000000000000000;
            14'h183c: o_data_a = 16'b1111110010101000;
            14'h183d: o_data_a = 16'b1111110000010000;
            14'h183e: o_data_a = 16'b0000000000000001;
            14'h183f: o_data_a = 16'b1111110111100000;
            14'h1840: o_data_a = 16'b1110001100001000;
            14'h1841: o_data_a = 16'b0000000000000000;
            14'h1842: o_data_a = 16'b1110110000010000;
            14'h1843: o_data_a = 16'b0000000000001101;
            14'h1844: o_data_a = 16'b1110001100001000;
            14'h1845: o_data_a = 16'b0110100110100010;
            14'h1846: o_data_a = 16'b1110110000010000;
            14'h1847: o_data_a = 16'b0000000000001110;
            14'h1848: o_data_a = 16'b1110001100001000;
            14'h1849: o_data_a = 16'b0001100001001101;
            14'h184a: o_data_a = 16'b1110110000010000;
            14'h184b: o_data_a = 16'b0000000001011111;
            14'h184c: o_data_a = 16'b1110101010000111;
            14'h184d: o_data_a = 16'b0000000000000000;
            14'h184e: o_data_a = 16'b1111110010101000;
            14'h184f: o_data_a = 16'b1111110000010000;
            14'h1850: o_data_a = 16'b0000000000000001;
            14'h1851: o_data_a = 16'b1111110111100000;
            14'h1852: o_data_a = 16'b1110110111100000;
            14'h1853: o_data_a = 16'b1110001100001000;
            14'h1854: o_data_a = 16'b0000000000000001;
            14'h1855: o_data_a = 16'b1111110000010000;
            14'h1856: o_data_a = 16'b0000000000000100;
            14'h1857: o_data_a = 16'b1110000010100000;
            14'h1858: o_data_a = 16'b1111110000010000;
            14'h1859: o_data_a = 16'b0000000000000000;
            14'h185a: o_data_a = 16'b1111110111101000;
            14'h185b: o_data_a = 16'b1110110010100000;
            14'h185c: o_data_a = 16'b1110001100001000;
            14'h185d: o_data_a = 16'b0000000000000000;
            14'h185e: o_data_a = 16'b1111110010100000;
            14'h185f: o_data_a = 16'b1111110001001000;
            14'h1860: o_data_a = 16'b0000000000000000;
            14'h1861: o_data_a = 16'b1111110010100000;
            14'h1862: o_data_a = 16'b1111110001001000;
            14'h1863: o_data_a = 16'b0000000000000000;
            14'h1864: o_data_a = 16'b1111110010101000;
            14'h1865: o_data_a = 16'b1111110000010000;
            14'h1866: o_data_a = 16'b0001100100000100;
            14'h1867: o_data_a = 16'b1110001100000101;
            14'h1868: o_data_a = 16'b0000000000000000;
            14'h1869: o_data_a = 16'b1110110000010000;
            14'h186a: o_data_a = 16'b0000000000001101;
            14'h186b: o_data_a = 16'b1110001100001000;
            14'h186c: o_data_a = 16'b0001011100111000;
            14'h186d: o_data_a = 16'b1110110000010000;
            14'h186e: o_data_a = 16'b0000000000001110;
            14'h186f: o_data_a = 16'b1110001100001000;
            14'h1870: o_data_a = 16'b0001100001110100;
            14'h1871: o_data_a = 16'b1110110000010000;
            14'h1872: o_data_a = 16'b0000000001011111;
            14'h1873: o_data_a = 16'b1110101010000111;
            14'h1874: o_data_a = 16'b0000000000000000;
            14'h1875: o_data_a = 16'b1111110010101000;
            14'h1876: o_data_a = 16'b1111110000010000;
            14'h1877: o_data_a = 16'b0000000000000001;
            14'h1878: o_data_a = 16'b1111110000100000;
            14'h1879: o_data_a = 16'b1110001100001000;
            14'h187a: o_data_a = 16'b0000000000000001;
            14'h187b: o_data_a = 16'b1111110000100000;
            14'h187c: o_data_a = 16'b1111110000010000;
            14'h187d: o_data_a = 16'b0000000000000000;
            14'h187e: o_data_a = 16'b1111110111101000;
            14'h187f: o_data_a = 16'b1110110010100000;
            14'h1880: o_data_a = 16'b1110001100001000;
            14'h1881: o_data_a = 16'b0000000000000001;
            14'h1882: o_data_a = 16'b1111110111100000;
            14'h1883: o_data_a = 16'b1111110000010000;
            14'h1884: o_data_a = 16'b0000000000000000;
            14'h1885: o_data_a = 16'b1111110111101000;
            14'h1886: o_data_a = 16'b1110110010100000;
            14'h1887: o_data_a = 16'b1110001100001000;
            14'h1888: o_data_a = 16'b0001100010001100;
            14'h1889: o_data_a = 16'b1110110000010000;
            14'h188a: o_data_a = 16'b0000000000000110;
            14'h188b: o_data_a = 16'b1110101010000111;
            14'h188c: o_data_a = 16'b0000000000000000;
            14'h188d: o_data_a = 16'b1111110010101000;
            14'h188e: o_data_a = 16'b1111110000010000;
            14'h188f: o_data_a = 16'b0000000000000001;
            14'h1890: o_data_a = 16'b1111110111100000;
            14'h1891: o_data_a = 16'b1110110111100000;
            14'h1892: o_data_a = 16'b1110110111100000;
            14'h1893: o_data_a = 16'b1110110111100000;
            14'h1894: o_data_a = 16'b1110001100001000;
            14'h1895: o_data_a = 16'b0000000000000001;
            14'h1896: o_data_a = 16'b1111110000010000;
            14'h1897: o_data_a = 16'b0000000000000100;
            14'h1898: o_data_a = 16'b1110000010100000;
            14'h1899: o_data_a = 16'b1111110000010000;
            14'h189a: o_data_a = 16'b0000000000000000;
            14'h189b: o_data_a = 16'b1111110111101000;
            14'h189c: o_data_a = 16'b1110110010100000;
            14'h189d: o_data_a = 16'b1110001100001000;
            14'h189e: o_data_a = 16'b0000000000000000;
            14'h189f: o_data_a = 16'b1111110010100000;
            14'h18a0: o_data_a = 16'b1111110001001000;
            14'h18a1: o_data_a = 16'b0000000000000000;
            14'h18a2: o_data_a = 16'b1111110010101000;
            14'h18a3: o_data_a = 16'b1111110000010000;
            14'h18a4: o_data_a = 16'b0001100010101000;
            14'h18a5: o_data_a = 16'b1110001100000101;
            14'h18a6: o_data_a = 16'b0001100100000010;
            14'h18a7: o_data_a = 16'b1110101010000111;
            14'h18a8: o_data_a = 16'b0000000000000001;
            14'h18a9: o_data_a = 16'b1111110000100000;
            14'h18aa: o_data_a = 16'b1111110000010000;
            14'h18ab: o_data_a = 16'b0000000000000000;
            14'h18ac: o_data_a = 16'b1111110111101000;
            14'h18ad: o_data_a = 16'b1110110010100000;
            14'h18ae: o_data_a = 16'b1110001100001000;
            14'h18af: o_data_a = 16'b0000000000000001;
            14'h18b0: o_data_a = 16'b1111110111100000;
            14'h18b1: o_data_a = 16'b1110110111100000;
            14'h18b2: o_data_a = 16'b1111110000010000;
            14'h18b3: o_data_a = 16'b0000000000000000;
            14'h18b4: o_data_a = 16'b1111110111101000;
            14'h18b5: o_data_a = 16'b1110110010100000;
            14'h18b6: o_data_a = 16'b1110001100001000;
            14'h18b7: o_data_a = 16'b0001100010111011;
            14'h18b8: o_data_a = 16'b1110110000010000;
            14'h18b9: o_data_a = 16'b0000000000000110;
            14'h18ba: o_data_a = 16'b1110101010000111;
            14'h18bb: o_data_a = 16'b0000000000000000;
            14'h18bc: o_data_a = 16'b1111110010101000;
            14'h18bd: o_data_a = 16'b1111110000010000;
            14'h18be: o_data_a = 16'b0001100011000010;
            14'h18bf: o_data_a = 16'b1110001100000101;
            14'h18c0: o_data_a = 16'b0001100011011110;
            14'h18c1: o_data_a = 16'b1110101010000111;
            14'h18c2: o_data_a = 16'b0000000000000001;
            14'h18c3: o_data_a = 16'b1111110000010000;
            14'h18c4: o_data_a = 16'b0000000000000011;
            14'h18c5: o_data_a = 16'b1110000010100000;
            14'h18c6: o_data_a = 16'b1111110000010000;
            14'h18c7: o_data_a = 16'b0000000000000000;
            14'h18c8: o_data_a = 16'b1111110111101000;
            14'h18c9: o_data_a = 16'b1110110010100000;
            14'h18ca: o_data_a = 16'b1110001100001000;
            14'h18cb: o_data_a = 16'b0000000000000001;
            14'h18cc: o_data_a = 16'b1110110000010000;
            14'h18cd: o_data_a = 16'b0000000000001101;
            14'h18ce: o_data_a = 16'b1110001100001000;
            14'h18cf: o_data_a = 16'b0110010011001001;
            14'h18d0: o_data_a = 16'b1110110000010000;
            14'h18d1: o_data_a = 16'b0000000000001110;
            14'h18d2: o_data_a = 16'b1110001100001000;
            14'h18d3: o_data_a = 16'b0001100011010111;
            14'h18d4: o_data_a = 16'b1110110000010000;
            14'h18d5: o_data_a = 16'b0000000001011111;
            14'h18d6: o_data_a = 16'b1110101010000111;
            14'h18d7: o_data_a = 16'b0000000000000000;
            14'h18d8: o_data_a = 16'b1111110010101000;
            14'h18d9: o_data_a = 16'b1111110000010000;
            14'h18da: o_data_a = 16'b0000000000000101;
            14'h18db: o_data_a = 16'b1110001100001000;
            14'h18dc: o_data_a = 16'b0001100100000010;
            14'h18dd: o_data_a = 16'b1110101010000111;
            14'h18de: o_data_a = 16'b0000000000000001;
            14'h18df: o_data_a = 16'b1111110000010000;
            14'h18e0: o_data_a = 16'b0000000000000011;
            14'h18e1: o_data_a = 16'b1110000010100000;
            14'h18e2: o_data_a = 16'b1111110000010000;
            14'h18e3: o_data_a = 16'b0000000000000000;
            14'h18e4: o_data_a = 16'b1111110111101000;
            14'h18e5: o_data_a = 16'b1110110010100000;
            14'h18e6: o_data_a = 16'b1110001100001000;
            14'h18e7: o_data_a = 16'b0000000000000001;
            14'h18e8: o_data_a = 16'b1111110000100000;
            14'h18e9: o_data_a = 16'b1111110000010000;
            14'h18ea: o_data_a = 16'b0000000000000000;
            14'h18eb: o_data_a = 16'b1111110111101000;
            14'h18ec: o_data_a = 16'b1110110010100000;
            14'h18ed: o_data_a = 16'b1110001100001000;
            14'h18ee: o_data_a = 16'b0000000000000010;
            14'h18ef: o_data_a = 16'b1110110000010000;
            14'h18f0: o_data_a = 16'b0000000000001101;
            14'h18f1: o_data_a = 16'b1110001100001000;
            14'h18f2: o_data_a = 16'b0110010000111011;
            14'h18f3: o_data_a = 16'b1110110000010000;
            14'h18f4: o_data_a = 16'b0000000000001110;
            14'h18f5: o_data_a = 16'b1110001100001000;
            14'h18f6: o_data_a = 16'b0001100011111010;
            14'h18f7: o_data_a = 16'b1110110000010000;
            14'h18f8: o_data_a = 16'b0000000001011111;
            14'h18f9: o_data_a = 16'b1110101010000111;
            14'h18fa: o_data_a = 16'b0000000000000000;
            14'h18fb: o_data_a = 16'b1111110010101000;
            14'h18fc: o_data_a = 16'b1111110000010000;
            14'h18fd: o_data_a = 16'b0000000000000001;
            14'h18fe: o_data_a = 16'b1111110111100000;
            14'h18ff: o_data_a = 16'b1110110111100000;
            14'h1900: o_data_a = 16'b1110110111100000;
            14'h1901: o_data_a = 16'b1110001100001000;
            14'h1902: o_data_a = 16'b0001100001010100;
            14'h1903: o_data_a = 16'b1110101010000111;
            14'h1904: o_data_a = 16'b0000000000000001;
            14'h1905: o_data_a = 16'b1111110000010000;
            14'h1906: o_data_a = 16'b0000000000000011;
            14'h1907: o_data_a = 16'b1110000010100000;
            14'h1908: o_data_a = 16'b1111110000010000;
            14'h1909: o_data_a = 16'b0000000000000000;
            14'h190a: o_data_a = 16'b1111110111101000;
            14'h190b: o_data_a = 16'b1110110010100000;
            14'h190c: o_data_a = 16'b1110001100001000;
            14'h190d: o_data_a = 16'b0000000000110110;
            14'h190e: o_data_a = 16'b1110101010000111;
            14'h190f: o_data_a = 16'b0000000000000000;
            14'h1910: o_data_a = 16'b1111110000100000;
            14'h1911: o_data_a = 16'b1110101010001000;
            14'h1912: o_data_a = 16'b1110110111110000;
            14'h1913: o_data_a = 16'b1110101010001000;
            14'h1914: o_data_a = 16'b0000000000000000;
            14'h1915: o_data_a = 16'b1110011111001000;
            14'h1916: o_data_a = 16'b0000000000000010;
            14'h1917: o_data_a = 16'b1111110000100000;
            14'h1918: o_data_a = 16'b1111110000010000;
            14'h1919: o_data_a = 16'b0000000000000000;
            14'h191a: o_data_a = 16'b1111110111101000;
            14'h191b: o_data_a = 16'b1110110010100000;
            14'h191c: o_data_a = 16'b1110001100001000;
            14'h191d: o_data_a = 16'b0000000000000001;
            14'h191e: o_data_a = 16'b1110110000010000;
            14'h191f: o_data_a = 16'b0000000000001101;
            14'h1920: o_data_a = 16'b1110001100001000;
            14'h1921: o_data_a = 16'b0001011111110100;
            14'h1922: o_data_a = 16'b1110110000010000;
            14'h1923: o_data_a = 16'b0000000000001110;
            14'h1924: o_data_a = 16'b1110001100001000;
            14'h1925: o_data_a = 16'b0001100100101001;
            14'h1926: o_data_a = 16'b1110110000010000;
            14'h1927: o_data_a = 16'b0000000001011111;
            14'h1928: o_data_a = 16'b1110101010000111;
            14'h1929: o_data_a = 16'b0000000000000000;
            14'h192a: o_data_a = 16'b1111110010101000;
            14'h192b: o_data_a = 16'b1111110000010000;
            14'h192c: o_data_a = 16'b0000000000000001;
            14'h192d: o_data_a = 16'b1111110000100000;
            14'h192e: o_data_a = 16'b1110001100001000;
            14'h192f: o_data_a = 16'b0000000000000001;
            14'h1930: o_data_a = 16'b1111110000100000;
            14'h1931: o_data_a = 16'b1111110000010000;
            14'h1932: o_data_a = 16'b0000000000000000;
            14'h1933: o_data_a = 16'b1111110111101000;
            14'h1934: o_data_a = 16'b1110110010100000;
            14'h1935: o_data_a = 16'b1110001100001000;
            14'h1936: o_data_a = 16'b0000000000000001;
            14'h1937: o_data_a = 16'b1110110000010000;
            14'h1938: o_data_a = 16'b0000000000001101;
            14'h1939: o_data_a = 16'b1110001100001000;
            14'h193a: o_data_a = 16'b0110010100100001;
            14'h193b: o_data_a = 16'b1110110000010000;
            14'h193c: o_data_a = 16'b0000000000001110;
            14'h193d: o_data_a = 16'b1110001100001000;
            14'h193e: o_data_a = 16'b0001100101000010;
            14'h193f: o_data_a = 16'b1110110000010000;
            14'h1940: o_data_a = 16'b0000000001011111;
            14'h1941: o_data_a = 16'b1110101010000111;
            14'h1942: o_data_a = 16'b0000000000000000;
            14'h1943: o_data_a = 16'b1111110010101000;
            14'h1944: o_data_a = 16'b1111110000010000;
            14'h1945: o_data_a = 16'b0000000000000001;
            14'h1946: o_data_a = 16'b1111110111100000;
            14'h1947: o_data_a = 16'b1110001100001000;
            14'h1948: o_data_a = 16'b0000000000000001;
            14'h1949: o_data_a = 16'b1111110000100000;
            14'h194a: o_data_a = 16'b1111110000010000;
            14'h194b: o_data_a = 16'b0000000000000000;
            14'h194c: o_data_a = 16'b1111110111101000;
            14'h194d: o_data_a = 16'b1110110010100000;
            14'h194e: o_data_a = 16'b1110001100001000;
            14'h194f: o_data_a = 16'b0000000000000001;
            14'h1950: o_data_a = 16'b1110110000010000;
            14'h1951: o_data_a = 16'b0000000000001101;
            14'h1952: o_data_a = 16'b1110001100001000;
            14'h1953: o_data_a = 16'b0110001010100100;
            14'h1954: o_data_a = 16'b1110110000010000;
            14'h1955: o_data_a = 16'b0000000000001110;
            14'h1956: o_data_a = 16'b1110001100001000;
            14'h1957: o_data_a = 16'b0001100101011011;
            14'h1958: o_data_a = 16'b1110110000010000;
            14'h1959: o_data_a = 16'b0000000001011111;
            14'h195a: o_data_a = 16'b1110101010000111;
            14'h195b: o_data_a = 16'b0000000000000000;
            14'h195c: o_data_a = 16'b1111110010101000;
            14'h195d: o_data_a = 16'b1111110000010000;
            14'h195e: o_data_a = 16'b0000000000000101;
            14'h195f: o_data_a = 16'b1110001100001000;
            14'h1960: o_data_a = 16'b0000000000000001;
            14'h1961: o_data_a = 16'b1111110111100000;
            14'h1962: o_data_a = 16'b1111110000010000;
            14'h1963: o_data_a = 16'b0000000000000000;
            14'h1964: o_data_a = 16'b1111110111101000;
            14'h1965: o_data_a = 16'b1110110010100000;
            14'h1966: o_data_a = 16'b1110001100001000;
            14'h1967: o_data_a = 16'b0000000000110110;
            14'h1968: o_data_a = 16'b1110101010000111;
            14'h1969: o_data_a = 16'b0000000000000000;
            14'h196a: o_data_a = 16'b1111110111101000;
            14'h196b: o_data_a = 16'b1110110010100000;
            14'h196c: o_data_a = 16'b1110101010001000;
            14'h196d: o_data_a = 16'b0000000000010000;
            14'h196e: o_data_a = 16'b1110110000010000;
            14'h196f: o_data_a = 16'b0000000000000000;
            14'h1970: o_data_a = 16'b1111110111101000;
            14'h1971: o_data_a = 16'b1110110010100000;
            14'h1972: o_data_a = 16'b1110001100001000;
            14'h1973: o_data_a = 16'b0000000000000001;
            14'h1974: o_data_a = 16'b1110110000010000;
            14'h1975: o_data_a = 16'b0000000000001101;
            14'h1976: o_data_a = 16'b1110001100001000;
            14'h1977: o_data_a = 16'b0001011010110000;
            14'h1978: o_data_a = 16'b1110110000010000;
            14'h1979: o_data_a = 16'b0000000000001110;
            14'h197a: o_data_a = 16'b1110001100001000;
            14'h197b: o_data_a = 16'b0001100101111111;
            14'h197c: o_data_a = 16'b1110110000010000;
            14'h197d: o_data_a = 16'b0000000001011111;
            14'h197e: o_data_a = 16'b1110101010000111;
            14'h197f: o_data_a = 16'b0000000000000000;
            14'h1980: o_data_a = 16'b1111110010101000;
            14'h1981: o_data_a = 16'b1111110000010000;
            14'h1982: o_data_a = 16'b0000000000010001;
            14'h1983: o_data_a = 16'b1110001100001000;
            14'h1984: o_data_a = 16'b0000000000010000;
            14'h1985: o_data_a = 16'b1110110000010000;
            14'h1986: o_data_a = 16'b0000000000000000;
            14'h1987: o_data_a = 16'b1111110111101000;
            14'h1988: o_data_a = 16'b1110110010100000;
            14'h1989: o_data_a = 16'b1110001100001000;
            14'h198a: o_data_a = 16'b0000000000000001;
            14'h198b: o_data_a = 16'b1110110000010000;
            14'h198c: o_data_a = 16'b0000000000001101;
            14'h198d: o_data_a = 16'b1110001100001000;
            14'h198e: o_data_a = 16'b0001011010110000;
            14'h198f: o_data_a = 16'b1110110000010000;
            14'h1990: o_data_a = 16'b0000000000001110;
            14'h1991: o_data_a = 16'b1110001100001000;
            14'h1992: o_data_a = 16'b0001100110010110;
            14'h1993: o_data_a = 16'b1110110000010000;
            14'h1994: o_data_a = 16'b0000000001011111;
            14'h1995: o_data_a = 16'b1110101010000111;
            14'h1996: o_data_a = 16'b0000000000000000;
            14'h1997: o_data_a = 16'b1111110010101000;
            14'h1998: o_data_a = 16'b1111110000010000;
            14'h1999: o_data_a = 16'b0000000000010010;
            14'h199a: o_data_a = 16'b1110001100001000;
            14'h199b: o_data_a = 16'b0000000000000000;
            14'h199c: o_data_a = 16'b1111110111001000;
            14'h199d: o_data_a = 16'b1111110010100000;
            14'h199e: o_data_a = 16'b1110101010001000;
            14'h199f: o_data_a = 16'b0000000000010010;
            14'h19a0: o_data_a = 16'b1111110000010000;
            14'h19a1: o_data_a = 16'b0000000000000000;
            14'h19a2: o_data_a = 16'b1111110111101000;
            14'h19a3: o_data_a = 16'b1110110010100000;
            14'h19a4: o_data_a = 16'b1110001100001000;
            14'h19a5: o_data_a = 16'b0000000000000000;
            14'h19a6: o_data_a = 16'b1111110010101000;
            14'h19a7: o_data_a = 16'b1111110000010000;
            14'h19a8: o_data_a = 16'b1110110010100000;
            14'h19a9: o_data_a = 16'b1111000010001000;
            14'h19aa: o_data_a = 16'b0000000000000000;
            14'h19ab: o_data_a = 16'b1111110111001000;
            14'h19ac: o_data_a = 16'b1111110010100000;
            14'h19ad: o_data_a = 16'b1110111111001000;
            14'h19ae: o_data_a = 16'b0000000000000000;
            14'h19af: o_data_a = 16'b1111110010101000;
            14'h19b0: o_data_a = 16'b1111110000010000;
            14'h19b1: o_data_a = 16'b0000000000000101;
            14'h19b2: o_data_a = 16'b1110001100001000;
            14'h19b3: o_data_a = 16'b0000000000000000;
            14'h19b4: o_data_a = 16'b1111110010101000;
            14'h19b5: o_data_a = 16'b1111110000010000;
            14'h19b6: o_data_a = 16'b0000000000000100;
            14'h19b7: o_data_a = 16'b1110001100001000;
            14'h19b8: o_data_a = 16'b0000000000000101;
            14'h19b9: o_data_a = 16'b1111110000010000;
            14'h19ba: o_data_a = 16'b0000000000000000;
            14'h19bb: o_data_a = 16'b1111110111101000;
            14'h19bc: o_data_a = 16'b1110110010100000;
            14'h19bd: o_data_a = 16'b1110001100001000;
            14'h19be: o_data_a = 16'b0000000000000000;
            14'h19bf: o_data_a = 16'b1111110010101000;
            14'h19c0: o_data_a = 16'b1111110000010000;
            14'h19c1: o_data_a = 16'b0000000000000100;
            14'h19c2: o_data_a = 16'b1111110000100000;
            14'h19c3: o_data_a = 16'b1110001100001000;
            14'h19c4: o_data_a = 16'b0000000000000001;
            14'h19c5: o_data_a = 16'b1111110000100000;
            14'h19c6: o_data_a = 16'b1111110000010000;
            14'h19c7: o_data_a = 16'b0000000000000000;
            14'h19c8: o_data_a = 16'b1111110111101000;
            14'h19c9: o_data_a = 16'b1110110010100000;
            14'h19ca: o_data_a = 16'b1110001100001000;
            14'h19cb: o_data_a = 16'b0000000000001111;
            14'h19cc: o_data_a = 16'b1110110000010000;
            14'h19cd: o_data_a = 16'b0000000000000000;
            14'h19ce: o_data_a = 16'b1111110111101000;
            14'h19cf: o_data_a = 16'b1110110010100000;
            14'h19d0: o_data_a = 16'b1110001100001000;
            14'h19d1: o_data_a = 16'b0001100111010101;
            14'h19d2: o_data_a = 16'b1110110000010000;
            14'h19d3: o_data_a = 16'b0000000000100110;
            14'h19d4: o_data_a = 16'b1110101010000111;
            14'h19d5: o_data_a = 16'b0000000000000000;
            14'h19d6: o_data_a = 16'b1111110010100000;
            14'h19d7: o_data_a = 16'b1111110001001000;
            14'h19d8: o_data_a = 16'b0000000000000000;
            14'h19d9: o_data_a = 16'b1111110010101000;
            14'h19da: o_data_a = 16'b1111110000010000;
            14'h19db: o_data_a = 16'b0001101001110000;
            14'h19dc: o_data_a = 16'b1110001100000101;
            14'h19dd: o_data_a = 16'b0000000000000001;
            14'h19de: o_data_a = 16'b1111110000100000;
            14'h19df: o_data_a = 16'b1111110000010000;
            14'h19e0: o_data_a = 16'b0000000000000000;
            14'h19e1: o_data_a = 16'b1111110111101000;
            14'h19e2: o_data_a = 16'b1110110010100000;
            14'h19e3: o_data_a = 16'b1110001100001000;
            14'h19e4: o_data_a = 16'b0000000000000000;
            14'h19e5: o_data_a = 16'b1111110111001000;
            14'h19e6: o_data_a = 16'b1111110010100000;
            14'h19e7: o_data_a = 16'b1110111111001000;
            14'h19e8: o_data_a = 16'b0000000000000000;
            14'h19e9: o_data_a = 16'b1111110010101000;
            14'h19ea: o_data_a = 16'b1111110000010000;
            14'h19eb: o_data_a = 16'b1110110010100000;
            14'h19ec: o_data_a = 16'b1111000010001000;
            14'h19ed: o_data_a = 16'b0000000000000000;
            14'h19ee: o_data_a = 16'b1111110010101000;
            14'h19ef: o_data_a = 16'b1111110000010000;
            14'h19f0: o_data_a = 16'b0000000000000001;
            14'h19f1: o_data_a = 16'b1111110000100000;
            14'h19f2: o_data_a = 16'b1110001100001000;
            14'h19f3: o_data_a = 16'b0000000000000001;
            14'h19f4: o_data_a = 16'b1111110000100000;
            14'h19f5: o_data_a = 16'b1111110000010000;
            14'h19f6: o_data_a = 16'b0000000000000000;
            14'h19f7: o_data_a = 16'b1111110111101000;
            14'h19f8: o_data_a = 16'b1110110010100000;
            14'h19f9: o_data_a = 16'b1110001100001000;
            14'h19fa: o_data_a = 16'b0000000000010010;
            14'h19fb: o_data_a = 16'b1111110000010000;
            14'h19fc: o_data_a = 16'b0000000000000000;
            14'h19fd: o_data_a = 16'b1111110111101000;
            14'h19fe: o_data_a = 16'b1110110010100000;
            14'h19ff: o_data_a = 16'b1110001100001000;
            14'h1a00: o_data_a = 16'b0000000000000000;
            14'h1a01: o_data_a = 16'b1111110010101000;
            14'h1a02: o_data_a = 16'b1111110000010000;
            14'h1a03: o_data_a = 16'b1110110010100000;
            14'h1a04: o_data_a = 16'b1111000010001000;
            14'h1a05: o_data_a = 16'b0000000000000001;
            14'h1a06: o_data_a = 16'b1111110000100000;
            14'h1a07: o_data_a = 16'b1111110000010000;
            14'h1a08: o_data_a = 16'b0000000000000000;
            14'h1a09: o_data_a = 16'b1111110111101000;
            14'h1a0a: o_data_a = 16'b1110110010100000;
            14'h1a0b: o_data_a = 16'b1110001100001000;
            14'h1a0c: o_data_a = 16'b0000000000000000;
            14'h1a0d: o_data_a = 16'b1111110111001000;
            14'h1a0e: o_data_a = 16'b1111110010100000;
            14'h1a0f: o_data_a = 16'b1110111111001000;
            14'h1a10: o_data_a = 16'b0000000000000000;
            14'h1a11: o_data_a = 16'b1111110010101000;
            14'h1a12: o_data_a = 16'b1111110000010000;
            14'h1a13: o_data_a = 16'b1110110010100000;
            14'h1a14: o_data_a = 16'b1111000111001000;
            14'h1a15: o_data_a = 16'b0000000000010010;
            14'h1a16: o_data_a = 16'b1111110000010000;
            14'h1a17: o_data_a = 16'b0000000000000000;
            14'h1a18: o_data_a = 16'b1111110111101000;
            14'h1a19: o_data_a = 16'b1110110010100000;
            14'h1a1a: o_data_a = 16'b1110001100001000;
            14'h1a1b: o_data_a = 16'b0000000000000000;
            14'h1a1c: o_data_a = 16'b1111110010101000;
            14'h1a1d: o_data_a = 16'b1111110000010000;
            14'h1a1e: o_data_a = 16'b1110110010100000;
            14'h1a1f: o_data_a = 16'b1111000010001000;
            14'h1a20: o_data_a = 16'b0000000000000000;
            14'h1a21: o_data_a = 16'b1111110010101000;
            14'h1a22: o_data_a = 16'b1111110000010000;
            14'h1a23: o_data_a = 16'b0000000000000100;
            14'h1a24: o_data_a = 16'b1110001100001000;
            14'h1a25: o_data_a = 16'b0000000000000100;
            14'h1a26: o_data_a = 16'b1111110000100000;
            14'h1a27: o_data_a = 16'b1111110000010000;
            14'h1a28: o_data_a = 16'b0000000000000000;
            14'h1a29: o_data_a = 16'b1111110111101000;
            14'h1a2a: o_data_a = 16'b1110110010100000;
            14'h1a2b: o_data_a = 16'b1110001100001000;
            14'h1a2c: o_data_a = 16'b0000000000000001;
            14'h1a2d: o_data_a = 16'b1111110000100000;
            14'h1a2e: o_data_a = 16'b1111110000010000;
            14'h1a2f: o_data_a = 16'b0000000000000000;
            14'h1a30: o_data_a = 16'b1111110111101000;
            14'h1a31: o_data_a = 16'b1110110010100000;
            14'h1a32: o_data_a = 16'b1110001100001000;
            14'h1a33: o_data_a = 16'b0000000000000000;
            14'h1a34: o_data_a = 16'b1111110111001000;
            14'h1a35: o_data_a = 16'b1111110010100000;
            14'h1a36: o_data_a = 16'b1110111111001000;
            14'h1a37: o_data_a = 16'b0000000000000000;
            14'h1a38: o_data_a = 16'b1111110010101000;
            14'h1a39: o_data_a = 16'b1111110000010000;
            14'h1a3a: o_data_a = 16'b1110110010100000;
            14'h1a3b: o_data_a = 16'b1111000111001000;
            14'h1a3c: o_data_a = 16'b0000000000010010;
            14'h1a3d: o_data_a = 16'b1111110000010000;
            14'h1a3e: o_data_a = 16'b0000000000000000;
            14'h1a3f: o_data_a = 16'b1111110111101000;
            14'h1a40: o_data_a = 16'b1110110010100000;
            14'h1a41: o_data_a = 16'b1110001100001000;
            14'h1a42: o_data_a = 16'b0000000000000000;
            14'h1a43: o_data_a = 16'b1111110010101000;
            14'h1a44: o_data_a = 16'b1111110000010000;
            14'h1a45: o_data_a = 16'b1110110010100000;
            14'h1a46: o_data_a = 16'b1111000010001000;
            14'h1a47: o_data_a = 16'b0000000000000000;
            14'h1a48: o_data_a = 16'b1111110010101000;
            14'h1a49: o_data_a = 16'b1111110000010000;
            14'h1a4a: o_data_a = 16'b0000000000000100;
            14'h1a4b: o_data_a = 16'b1110001100001000;
            14'h1a4c: o_data_a = 16'b0000000000000100;
            14'h1a4d: o_data_a = 16'b1111110000100000;
            14'h1a4e: o_data_a = 16'b1111110000010000;
            14'h1a4f: o_data_a = 16'b0000000000000000;
            14'h1a50: o_data_a = 16'b1111110111101000;
            14'h1a51: o_data_a = 16'b1110110010100000;
            14'h1a52: o_data_a = 16'b1110001100001000;
            14'h1a53: o_data_a = 16'b0000000000000000;
            14'h1a54: o_data_a = 16'b1111110010101000;
            14'h1a55: o_data_a = 16'b1111110000010000;
            14'h1a56: o_data_a = 16'b1110110010100000;
            14'h1a57: o_data_a = 16'b1111000010001000;
            14'h1a58: o_data_a = 16'b0000000000000000;
            14'h1a59: o_data_a = 16'b1111110010101000;
            14'h1a5a: o_data_a = 16'b1111110000010000;
            14'h1a5b: o_data_a = 16'b0000000000000101;
            14'h1a5c: o_data_a = 16'b1110001100001000;
            14'h1a5d: o_data_a = 16'b0000000000000000;
            14'h1a5e: o_data_a = 16'b1111110010101000;
            14'h1a5f: o_data_a = 16'b1111110000010000;
            14'h1a60: o_data_a = 16'b0000000000000100;
            14'h1a61: o_data_a = 16'b1110001100001000;
            14'h1a62: o_data_a = 16'b0000000000000101;
            14'h1a63: o_data_a = 16'b1111110000010000;
            14'h1a64: o_data_a = 16'b0000000000000000;
            14'h1a65: o_data_a = 16'b1111110111101000;
            14'h1a66: o_data_a = 16'b1110110010100000;
            14'h1a67: o_data_a = 16'b1110001100001000;
            14'h1a68: o_data_a = 16'b0000000000000000;
            14'h1a69: o_data_a = 16'b1111110010101000;
            14'h1a6a: o_data_a = 16'b1111110000010000;
            14'h1a6b: o_data_a = 16'b0000000000000100;
            14'h1a6c: o_data_a = 16'b1111110000100000;
            14'h1a6d: o_data_a = 16'b1110001100001000;
            14'h1a6e: o_data_a = 16'b0001100111000100;
            14'h1a6f: o_data_a = 16'b1110101010000111;
            14'h1a70: o_data_a = 16'b0000000000000000;
            14'h1a71: o_data_a = 16'b1111110111001000;
            14'h1a72: o_data_a = 16'b1111110010100000;
            14'h1a73: o_data_a = 16'b1110101010001000;
            14'h1a74: o_data_a = 16'b0000000000110110;
            14'h1a75: o_data_a = 16'b1110101010000111;
            14'h1a76: o_data_a = 16'b0000000000000010;
            14'h1a77: o_data_a = 16'b1111110000100000;
            14'h1a78: o_data_a = 16'b1111110000010000;
            14'h1a79: o_data_a = 16'b0000000000000000;
            14'h1a7a: o_data_a = 16'b1111110111101000;
            14'h1a7b: o_data_a = 16'b1110110010100000;
            14'h1a7c: o_data_a = 16'b1110001100001000;
            14'h1a7d: o_data_a = 16'b0000000000000000;
            14'h1a7e: o_data_a = 16'b1111110111001000;
            14'h1a7f: o_data_a = 16'b1111110010100000;
            14'h1a80: o_data_a = 16'b1110101010001000;
            14'h1a81: o_data_a = 16'b0001101010000101;
            14'h1a82: o_data_a = 16'b1110110000010000;
            14'h1a83: o_data_a = 16'b0000000000100110;
            14'h1a84: o_data_a = 16'b1110101010000111;
            14'h1a85: o_data_a = 16'b0000000000000000;
            14'h1a86: o_data_a = 16'b1111110010101000;
            14'h1a87: o_data_a = 16'b1111110000010000;
            14'h1a88: o_data_a = 16'b0001101010001100;
            14'h1a89: o_data_a = 16'b1110001100000101;
            14'h1a8a: o_data_a = 16'b0001101010011101;
            14'h1a8b: o_data_a = 16'b1110101010000111;
            14'h1a8c: o_data_a = 16'b0000000000000010;
            14'h1a8d: o_data_a = 16'b1111110000100000;
            14'h1a8e: o_data_a = 16'b1111110000010000;
            14'h1a8f: o_data_a = 16'b0000000000000000;
            14'h1a90: o_data_a = 16'b1111110111101000;
            14'h1a91: o_data_a = 16'b1110110010100000;
            14'h1a92: o_data_a = 16'b1110001100001000;
            14'h1a93: o_data_a = 16'b0000000000000000;
            14'h1a94: o_data_a = 16'b1111110010100000;
            14'h1a95: o_data_a = 16'b1111110001010000;
            14'h1a96: o_data_a = 16'b1110011111001000;
            14'h1a97: o_data_a = 16'b0000000000000000;
            14'h1a98: o_data_a = 16'b1111110010101000;
            14'h1a99: o_data_a = 16'b1111110000010000;
            14'h1a9a: o_data_a = 16'b0000000000000010;
            14'h1a9b: o_data_a = 16'b1111110000100000;
            14'h1a9c: o_data_a = 16'b1110001100001000;
            14'h1a9d: o_data_a = 16'b0000000000000010;
            14'h1a9e: o_data_a = 16'b1111110000100000;
            14'h1a9f: o_data_a = 16'b1111110000010000;
            14'h1aa0: o_data_a = 16'b0000000000000000;
            14'h1aa1: o_data_a = 16'b1111110111101000;
            14'h1aa2: o_data_a = 16'b1110110010100000;
            14'h1aa3: o_data_a = 16'b1110001100001000;
            14'h1aa4: o_data_a = 16'b0000000000110110;
            14'h1aa5: o_data_a = 16'b1110101010000111;
            14'h1aa6: o_data_a = 16'b0000000000000101;
            14'h1aa7: o_data_a = 16'b1110110000010000;
            14'h1aa8: o_data_a = 16'b1110001110010000;
            14'h1aa9: o_data_a = 16'b0000000000000000;
            14'h1aaa: o_data_a = 16'b1111110111101000;
            14'h1aab: o_data_a = 16'b1110110010100000;
            14'h1aac: o_data_a = 16'b1110101010001000;
            14'h1aad: o_data_a = 16'b0001101010101000;
            14'h1aae: o_data_a = 16'b1110001100000001;
            14'h1aaf: o_data_a = 16'b0000000000000010;
            14'h1ab0: o_data_a = 16'b1111110000100000;
            14'h1ab1: o_data_a = 16'b1111110000010000;
            14'h1ab2: o_data_a = 16'b0000000000000000;
            14'h1ab3: o_data_a = 16'b1111110111101000;
            14'h1ab4: o_data_a = 16'b1110110010100000;
            14'h1ab5: o_data_a = 16'b1110001100001000;
            14'h1ab6: o_data_a = 16'b0000000000000000;
            14'h1ab7: o_data_a = 16'b1111110111001000;
            14'h1ab8: o_data_a = 16'b1111110010100000;
            14'h1ab9: o_data_a = 16'b1110101010001000;
            14'h1aba: o_data_a = 16'b0001101010111110;
            14'h1abb: o_data_a = 16'b1110110000010000;
            14'h1abc: o_data_a = 16'b0000000000100110;
            14'h1abd: o_data_a = 16'b1110101010000111;
            14'h1abe: o_data_a = 16'b0000000000000010;
            14'h1abf: o_data_a = 16'b1111110111100000;
            14'h1ac0: o_data_a = 16'b1111110000010000;
            14'h1ac1: o_data_a = 16'b0000000000000000;
            14'h1ac2: o_data_a = 16'b1111110111101000;
            14'h1ac3: o_data_a = 16'b1110110010100000;
            14'h1ac4: o_data_a = 16'b1110001100001000;
            14'h1ac5: o_data_a = 16'b0000000000000000;
            14'h1ac6: o_data_a = 16'b1111110111001000;
            14'h1ac7: o_data_a = 16'b1111110010100000;
            14'h1ac8: o_data_a = 16'b1110101010001000;
            14'h1ac9: o_data_a = 16'b0001101011001101;
            14'h1aca: o_data_a = 16'b1110110000010000;
            14'h1acb: o_data_a = 16'b0000000000010110;
            14'h1acc: o_data_a = 16'b1110101010000111;
            14'h1acd: o_data_a = 16'b0000000000000000;
            14'h1ace: o_data_a = 16'b1111110010101000;
            14'h1acf: o_data_a = 16'b1111110000010000;
            14'h1ad0: o_data_a = 16'b1110110010100000;
            14'h1ad1: o_data_a = 16'b1111000000001000;
            14'h1ad2: o_data_a = 16'b0000000000000010;
            14'h1ad3: o_data_a = 16'b1111110000100000;
            14'h1ad4: o_data_a = 16'b1111110000010000;
            14'h1ad5: o_data_a = 16'b0000000000000000;
            14'h1ad6: o_data_a = 16'b1111110111101000;
            14'h1ad7: o_data_a = 16'b1110110010100000;
            14'h1ad8: o_data_a = 16'b1110001100001000;
            14'h1ad9: o_data_a = 16'b0000000000000000;
            14'h1ada: o_data_a = 16'b1111110111001000;
            14'h1adb: o_data_a = 16'b1111110010100000;
            14'h1adc: o_data_a = 16'b1110101010001000;
            14'h1add: o_data_a = 16'b0001101011100001;
            14'h1ade: o_data_a = 16'b1110110000010000;
            14'h1adf: o_data_a = 16'b0000000000010110;
            14'h1ae0: o_data_a = 16'b1110101010000111;
            14'h1ae1: o_data_a = 16'b0000000000000010;
            14'h1ae2: o_data_a = 16'b1111110111100000;
            14'h1ae3: o_data_a = 16'b1111110000010000;
            14'h1ae4: o_data_a = 16'b0000000000000000;
            14'h1ae5: o_data_a = 16'b1111110111101000;
            14'h1ae6: o_data_a = 16'b1110110010100000;
            14'h1ae7: o_data_a = 16'b1110001100001000;
            14'h1ae8: o_data_a = 16'b0000000000000000;
            14'h1ae9: o_data_a = 16'b1111110111001000;
            14'h1aea: o_data_a = 16'b1111110010100000;
            14'h1aeb: o_data_a = 16'b1110101010001000;
            14'h1aec: o_data_a = 16'b0001101011110000;
            14'h1aed: o_data_a = 16'b1110110000010000;
            14'h1aee: o_data_a = 16'b0000000000100110;
            14'h1aef: o_data_a = 16'b1110101010000111;
            14'h1af0: o_data_a = 16'b0000000000000000;
            14'h1af1: o_data_a = 16'b1111110010101000;
            14'h1af2: o_data_a = 16'b1111110000010000;
            14'h1af3: o_data_a = 16'b1110110010100000;
            14'h1af4: o_data_a = 16'b1111000000001000;
            14'h1af5: o_data_a = 16'b0000000000000000;
            14'h1af6: o_data_a = 16'b1111110010101000;
            14'h1af7: o_data_a = 16'b1111110000010000;
            14'h1af8: o_data_a = 16'b1110110010100000;
            14'h1af9: o_data_a = 16'b1111010101001000;
            14'h1afa: o_data_a = 16'b0000000000000000;
            14'h1afb: o_data_a = 16'b1111110010101000;
            14'h1afc: o_data_a = 16'b1111110000010000;
            14'h1afd: o_data_a = 16'b0000000000000001;
            14'h1afe: o_data_a = 16'b1111110111100000;
            14'h1aff: o_data_a = 16'b1110110111100000;
            14'h1b00: o_data_a = 16'b1110110111100000;
            14'h1b01: o_data_a = 16'b1110110111100000;
            14'h1b02: o_data_a = 16'b1110001100001000;
            14'h1b03: o_data_a = 16'b0000000000000010;
            14'h1b04: o_data_a = 16'b1111110000100000;
            14'h1b05: o_data_a = 16'b1111110000010000;
            14'h1b06: o_data_a = 16'b0000000000000000;
            14'h1b07: o_data_a = 16'b1111110111101000;
            14'h1b08: o_data_a = 16'b1110110010100000;
            14'h1b09: o_data_a = 16'b1110001100001000;
            14'h1b0a: o_data_a = 16'b0000000000000001;
            14'h1b0b: o_data_a = 16'b1110110000010000;
            14'h1b0c: o_data_a = 16'b0000000000001101;
            14'h1b0d: o_data_a = 16'b1110001100001000;
            14'h1b0e: o_data_a = 16'b0001101001110110;
            14'h1b0f: o_data_a = 16'b1110110000010000;
            14'h1b10: o_data_a = 16'b0000000000001110;
            14'h1b11: o_data_a = 16'b1110001100001000;
            14'h1b12: o_data_a = 16'b0001101100010110;
            14'h1b13: o_data_a = 16'b1110110000010000;
            14'h1b14: o_data_a = 16'b0000000001011111;
            14'h1b15: o_data_a = 16'b1110101010000111;
            14'h1b16: o_data_a = 16'b0000000000000000;
            14'h1b17: o_data_a = 16'b1111110010101000;
            14'h1b18: o_data_a = 16'b1111110000010000;
            14'h1b19: o_data_a = 16'b0000000000000010;
            14'h1b1a: o_data_a = 16'b1111110000100000;
            14'h1b1b: o_data_a = 16'b1110001100001000;
            14'h1b1c: o_data_a = 16'b0000000000000010;
            14'h1b1d: o_data_a = 16'b1111110111100000;
            14'h1b1e: o_data_a = 16'b1111110000010000;
            14'h1b1f: o_data_a = 16'b0000000000000000;
            14'h1b20: o_data_a = 16'b1111110111101000;
            14'h1b21: o_data_a = 16'b1110110010100000;
            14'h1b22: o_data_a = 16'b1110001100001000;
            14'h1b23: o_data_a = 16'b0000000000000001;
            14'h1b24: o_data_a = 16'b1110110000010000;
            14'h1b25: o_data_a = 16'b0000000000001101;
            14'h1b26: o_data_a = 16'b1110001100001000;
            14'h1b27: o_data_a = 16'b0001101001110110;
            14'h1b28: o_data_a = 16'b1110110000010000;
            14'h1b29: o_data_a = 16'b0000000000001110;
            14'h1b2a: o_data_a = 16'b1110001100001000;
            14'h1b2b: o_data_a = 16'b0001101100101111;
            14'h1b2c: o_data_a = 16'b1110110000010000;
            14'h1b2d: o_data_a = 16'b0000000001011111;
            14'h1b2e: o_data_a = 16'b1110101010000111;
            14'h1b2f: o_data_a = 16'b0000000000000000;
            14'h1b30: o_data_a = 16'b1111110010101000;
            14'h1b31: o_data_a = 16'b1111110000010000;
            14'h1b32: o_data_a = 16'b0000000000000010;
            14'h1b33: o_data_a = 16'b1111110111100000;
            14'h1b34: o_data_a = 16'b1110001100001000;
            14'h1b35: o_data_a = 16'b0000000000000010;
            14'h1b36: o_data_a = 16'b1111110000100000;
            14'h1b37: o_data_a = 16'b1111110000010000;
            14'h1b38: o_data_a = 16'b0000000000000000;
            14'h1b39: o_data_a = 16'b1111110111101000;
            14'h1b3a: o_data_a = 16'b1110110010100000;
            14'h1b3b: o_data_a = 16'b1110001100001000;
            14'h1b3c: o_data_a = 16'b0000000000000010;
            14'h1b3d: o_data_a = 16'b1111110111100000;
            14'h1b3e: o_data_a = 16'b1111110000010000;
            14'h1b3f: o_data_a = 16'b0000000000000000;
            14'h1b40: o_data_a = 16'b1111110111101000;
            14'h1b41: o_data_a = 16'b1110110010100000;
            14'h1b42: o_data_a = 16'b1110001100001000;
            14'h1b43: o_data_a = 16'b0001101101000111;
            14'h1b44: o_data_a = 16'b1110110000010000;
            14'h1b45: o_data_a = 16'b0000000000100110;
            14'h1b46: o_data_a = 16'b1110101010000111;
            14'h1b47: o_data_a = 16'b0000000000000000;
            14'h1b48: o_data_a = 16'b1111110010101000;
            14'h1b49: o_data_a = 16'b1111110000010000;
            14'h1b4a: o_data_a = 16'b0001101101001110;
            14'h1b4b: o_data_a = 16'b1110001100000101;
            14'h1b4c: o_data_a = 16'b0001101101110101;
            14'h1b4d: o_data_a = 16'b1110101010000111;
            14'h1b4e: o_data_a = 16'b0000000000000010;
            14'h1b4f: o_data_a = 16'b1111110000100000;
            14'h1b50: o_data_a = 16'b1111110000010000;
            14'h1b51: o_data_a = 16'b0000000000000000;
            14'h1b52: o_data_a = 16'b1111110111101000;
            14'h1b53: o_data_a = 16'b1110110010100000;
            14'h1b54: o_data_a = 16'b1110001100001000;
            14'h1b55: o_data_a = 16'b0000000000000000;
            14'h1b56: o_data_a = 16'b1111110010101000;
            14'h1b57: o_data_a = 16'b1111110000010000;
            14'h1b58: o_data_a = 16'b0000000000000001;
            14'h1b59: o_data_a = 16'b1111110111100000;
            14'h1b5a: o_data_a = 16'b1110001100001000;
            14'h1b5b: o_data_a = 16'b0000000000000010;
            14'h1b5c: o_data_a = 16'b1111110111100000;
            14'h1b5d: o_data_a = 16'b1111110000010000;
            14'h1b5e: o_data_a = 16'b0000000000000000;
            14'h1b5f: o_data_a = 16'b1111110111101000;
            14'h1b60: o_data_a = 16'b1110110010100000;
            14'h1b61: o_data_a = 16'b1110001100001000;
            14'h1b62: o_data_a = 16'b0000000000000000;
            14'h1b63: o_data_a = 16'b1111110010101000;
            14'h1b64: o_data_a = 16'b1111110000010000;
            14'h1b65: o_data_a = 16'b0000000000000010;
            14'h1b66: o_data_a = 16'b1111110000100000;
            14'h1b67: o_data_a = 16'b1110001100001000;
            14'h1b68: o_data_a = 16'b0000000000000001;
            14'h1b69: o_data_a = 16'b1111110111100000;
            14'h1b6a: o_data_a = 16'b1111110000010000;
            14'h1b6b: o_data_a = 16'b0000000000000000;
            14'h1b6c: o_data_a = 16'b1111110111101000;
            14'h1b6d: o_data_a = 16'b1110110010100000;
            14'h1b6e: o_data_a = 16'b1110001100001000;
            14'h1b6f: o_data_a = 16'b0000000000000000;
            14'h1b70: o_data_a = 16'b1111110010101000;
            14'h1b71: o_data_a = 16'b1111110000010000;
            14'h1b72: o_data_a = 16'b0000000000000010;
            14'h1b73: o_data_a = 16'b1111110111100000;
            14'h1b74: o_data_a = 16'b1110001100001000;
            14'h1b75: o_data_a = 16'b0000000000000001;
            14'h1b76: o_data_a = 16'b1111110111100000;
            14'h1b77: o_data_a = 16'b1110110111100000;
            14'h1b78: o_data_a = 16'b1111110000010000;
            14'h1b79: o_data_a = 16'b0000000000000000;
            14'h1b7a: o_data_a = 16'b1111110111101000;
            14'h1b7b: o_data_a = 16'b1110110010100000;
            14'h1b7c: o_data_a = 16'b1110001100001000;
            14'h1b7d: o_data_a = 16'b0000000000000010;
            14'h1b7e: o_data_a = 16'b1111110111100000;
            14'h1b7f: o_data_a = 16'b1111110000010000;
            14'h1b80: o_data_a = 16'b0000000000000000;
            14'h1b81: o_data_a = 16'b1111110111101000;
            14'h1b82: o_data_a = 16'b1110110010100000;
            14'h1b83: o_data_a = 16'b1110001100001000;
            14'h1b84: o_data_a = 16'b0001101110001000;
            14'h1b85: o_data_a = 16'b1110110000010000;
            14'h1b86: o_data_a = 16'b0000000000100110;
            14'h1b87: o_data_a = 16'b1110101010000111;
            14'h1b88: o_data_a = 16'b0000000000000000;
            14'h1b89: o_data_a = 16'b1111110010100000;
            14'h1b8a: o_data_a = 16'b1111110001001000;
            14'h1b8b: o_data_a = 16'b0000000000000000;
            14'h1b8c: o_data_a = 16'b1111110010101000;
            14'h1b8d: o_data_a = 16'b1111110000010000;
            14'h1b8e: o_data_a = 16'b0001110001001101;
            14'h1b8f: o_data_a = 16'b1110001100000101;
            14'h1b90: o_data_a = 16'b0000000000000001;
            14'h1b91: o_data_a = 16'b1111110000010000;
            14'h1b92: o_data_a = 16'b0000000000000011;
            14'h1b93: o_data_a = 16'b1110000010100000;
            14'h1b94: o_data_a = 16'b1111110000010000;
            14'h1b95: o_data_a = 16'b0000000000000000;
            14'h1b96: o_data_a = 16'b1111110111101000;
            14'h1b97: o_data_a = 16'b1110110010100000;
            14'h1b98: o_data_a = 16'b1110001100001000;
            14'h1b99: o_data_a = 16'b0000000000010010;
            14'h1b9a: o_data_a = 16'b1111110000010000;
            14'h1b9b: o_data_a = 16'b0000000000000000;
            14'h1b9c: o_data_a = 16'b1111110111101000;
            14'h1b9d: o_data_a = 16'b1110110010100000;
            14'h1b9e: o_data_a = 16'b1110001100001000;
            14'h1b9f: o_data_a = 16'b0000000000000000;
            14'h1ba0: o_data_a = 16'b1111110010101000;
            14'h1ba1: o_data_a = 16'b1111110000010000;
            14'h1ba2: o_data_a = 16'b1110110010100000;
            14'h1ba3: o_data_a = 16'b1111000010001000;
            14'h1ba4: o_data_a = 16'b0000000000000000;
            14'h1ba5: o_data_a = 16'b1111110010101000;
            14'h1ba6: o_data_a = 16'b1111110000010000;
            14'h1ba7: o_data_a = 16'b0000000000000100;
            14'h1ba8: o_data_a = 16'b1110001100001000;
            14'h1ba9: o_data_a = 16'b0000000000000100;
            14'h1baa: o_data_a = 16'b1111110000100000;
            14'h1bab: o_data_a = 16'b1111110000010000;
            14'h1bac: o_data_a = 16'b0000000000000000;
            14'h1bad: o_data_a = 16'b1111110111101000;
            14'h1bae: o_data_a = 16'b1110110010100000;
            14'h1baf: o_data_a = 16'b1110001100001000;
            14'h1bb0: o_data_a = 16'b0000000000000010;
            14'h1bb1: o_data_a = 16'b1111110111100000;
            14'h1bb2: o_data_a = 16'b1111110000010000;
            14'h1bb3: o_data_a = 16'b0000000000000000;
            14'h1bb4: o_data_a = 16'b1111110111101000;
            14'h1bb5: o_data_a = 16'b1110110010100000;
            14'h1bb6: o_data_a = 16'b1110001100001000;
            14'h1bb7: o_data_a = 16'b0000000000000000;
            14'h1bb8: o_data_a = 16'b1111110010101000;
            14'h1bb9: o_data_a = 16'b1111110000010000;
            14'h1bba: o_data_a = 16'b1110110010100000;
            14'h1bbb: o_data_a = 16'b1111000000001000;
            14'h1bbc: o_data_a = 16'b0000000000000000;
            14'h1bbd: o_data_a = 16'b1111110111001000;
            14'h1bbe: o_data_a = 16'b1111110010100000;
            14'h1bbf: o_data_a = 16'b1110101010001000;
            14'h1bc0: o_data_a = 16'b0001101111000100;
            14'h1bc1: o_data_a = 16'b1110110000010000;
            14'h1bc2: o_data_a = 16'b0000000000010110;
            14'h1bc3: o_data_a = 16'b1110101010000111;
            14'h1bc4: o_data_a = 16'b0000000000000000;
            14'h1bc5: o_data_a = 16'b1111110010101000;
            14'h1bc6: o_data_a = 16'b1111110000010000;
            14'h1bc7: o_data_a = 16'b0001101111001011;
            14'h1bc8: o_data_a = 16'b1110001100000101;
            14'h1bc9: o_data_a = 16'b0001110000011000;
            14'h1bca: o_data_a = 16'b1110101010000111;
            14'h1bcb: o_data_a = 16'b0000000000000001;
            14'h1bcc: o_data_a = 16'b1111110000100000;
            14'h1bcd: o_data_a = 16'b1111110000010000;
            14'h1bce: o_data_a = 16'b0000000000000000;
            14'h1bcf: o_data_a = 16'b1111110111101000;
            14'h1bd0: o_data_a = 16'b1110110010100000;
            14'h1bd1: o_data_a = 16'b1110001100001000;
            14'h1bd2: o_data_a = 16'b0000000000000010;
            14'h1bd3: o_data_a = 16'b1111110000100000;
            14'h1bd4: o_data_a = 16'b1111110000010000;
            14'h1bd5: o_data_a = 16'b0000000000000000;
            14'h1bd6: o_data_a = 16'b1111110111101000;
            14'h1bd7: o_data_a = 16'b1110110010100000;
            14'h1bd8: o_data_a = 16'b1110001100001000;
            14'h1bd9: o_data_a = 16'b0000000000000000;
            14'h1bda: o_data_a = 16'b1111110010101000;
            14'h1bdb: o_data_a = 16'b1111110000010000;
            14'h1bdc: o_data_a = 16'b1110110010100000;
            14'h1bdd: o_data_a = 16'b1111000010001000;
            14'h1bde: o_data_a = 16'b0000000000000000;
            14'h1bdf: o_data_a = 16'b1111110010101000;
            14'h1be0: o_data_a = 16'b1111110000010000;
            14'h1be1: o_data_a = 16'b0000000000000001;
            14'h1be2: o_data_a = 16'b1111110000100000;
            14'h1be3: o_data_a = 16'b1110001100001000;
            14'h1be4: o_data_a = 16'b0000000000000001;
            14'h1be5: o_data_a = 16'b1111110111100000;
            14'h1be6: o_data_a = 16'b1110110111100000;
            14'h1be7: o_data_a = 16'b1111110000010000;
            14'h1be8: o_data_a = 16'b0000000000000000;
            14'h1be9: o_data_a = 16'b1111110111101000;
            14'h1bea: o_data_a = 16'b1110110010100000;
            14'h1beb: o_data_a = 16'b1110001100001000;
            14'h1bec: o_data_a = 16'b0000000000000001;
            14'h1bed: o_data_a = 16'b1111110000010000;
            14'h1bee: o_data_a = 16'b0000000000000011;
            14'h1bef: o_data_a = 16'b1110000010100000;
            14'h1bf0: o_data_a = 16'b1111110000010000;
            14'h1bf1: o_data_a = 16'b0000000000000000;
            14'h1bf2: o_data_a = 16'b1111110111101000;
            14'h1bf3: o_data_a = 16'b1110110010100000;
            14'h1bf4: o_data_a = 16'b1110001100001000;
            14'h1bf5: o_data_a = 16'b0000000000010010;
            14'h1bf6: o_data_a = 16'b1111110000010000;
            14'h1bf7: o_data_a = 16'b0000000000000000;
            14'h1bf8: o_data_a = 16'b1111110111101000;
            14'h1bf9: o_data_a = 16'b1110110010100000;
            14'h1bfa: o_data_a = 16'b1110001100001000;
            14'h1bfb: o_data_a = 16'b0000000000000000;
            14'h1bfc: o_data_a = 16'b1111110010101000;
            14'h1bfd: o_data_a = 16'b1111110000010000;
            14'h1bfe: o_data_a = 16'b1110110010100000;
            14'h1bff: o_data_a = 16'b1111000010001000;
            14'h1c00: o_data_a = 16'b0000000000000000;
            14'h1c01: o_data_a = 16'b1111110010101000;
            14'h1c02: o_data_a = 16'b1111110000010000;
            14'h1c03: o_data_a = 16'b0000000000000100;
            14'h1c04: o_data_a = 16'b1110001100001000;
            14'h1c05: o_data_a = 16'b0000000000000100;
            14'h1c06: o_data_a = 16'b1111110000100000;
            14'h1c07: o_data_a = 16'b1111110000010000;
            14'h1c08: o_data_a = 16'b0000000000000000;
            14'h1c09: o_data_a = 16'b1111110111101000;
            14'h1c0a: o_data_a = 16'b1110110010100000;
            14'h1c0b: o_data_a = 16'b1110001100001000;
            14'h1c0c: o_data_a = 16'b0000000000000000;
            14'h1c0d: o_data_a = 16'b1111110010101000;
            14'h1c0e: o_data_a = 16'b1111110000010000;
            14'h1c0f: o_data_a = 16'b1110110010100000;
            14'h1c10: o_data_a = 16'b1111000010001000;
            14'h1c11: o_data_a = 16'b0000000000000000;
            14'h1c12: o_data_a = 16'b1111110010101000;
            14'h1c13: o_data_a = 16'b1111110000010000;
            14'h1c14: o_data_a = 16'b0000000000000001;
            14'h1c15: o_data_a = 16'b1111110111100000;
            14'h1c16: o_data_a = 16'b1110110111100000;
            14'h1c17: o_data_a = 16'b1110001100001000;
            14'h1c18: o_data_a = 16'b0000000000000010;
            14'h1c19: o_data_a = 16'b1111110000100000;
            14'h1c1a: o_data_a = 16'b1111110000010000;
            14'h1c1b: o_data_a = 16'b0000000000000000;
            14'h1c1c: o_data_a = 16'b1111110111101000;
            14'h1c1d: o_data_a = 16'b1110110010100000;
            14'h1c1e: o_data_a = 16'b1110001100001000;
            14'h1c1f: o_data_a = 16'b0000000000000010;
            14'h1c20: o_data_a = 16'b1111110000100000;
            14'h1c21: o_data_a = 16'b1111110000010000;
            14'h1c22: o_data_a = 16'b0000000000000000;
            14'h1c23: o_data_a = 16'b1111110111101000;
            14'h1c24: o_data_a = 16'b1110110010100000;
            14'h1c25: o_data_a = 16'b1110001100001000;
            14'h1c26: o_data_a = 16'b0000000000000000;
            14'h1c27: o_data_a = 16'b1111110010101000;
            14'h1c28: o_data_a = 16'b1111110000010000;
            14'h1c29: o_data_a = 16'b1110110010100000;
            14'h1c2a: o_data_a = 16'b1111000010001000;
            14'h1c2b: o_data_a = 16'b0000000000000000;
            14'h1c2c: o_data_a = 16'b1111110010101000;
            14'h1c2d: o_data_a = 16'b1111110000010000;
            14'h1c2e: o_data_a = 16'b0000000000000010;
            14'h1c2f: o_data_a = 16'b1111110000100000;
            14'h1c30: o_data_a = 16'b1110001100001000;
            14'h1c31: o_data_a = 16'b0000000000000001;
            14'h1c32: o_data_a = 16'b1111110000010000;
            14'h1c33: o_data_a = 16'b0000000000000011;
            14'h1c34: o_data_a = 16'b1110000010100000;
            14'h1c35: o_data_a = 16'b1111110000010000;
            14'h1c36: o_data_a = 16'b0000000000000000;
            14'h1c37: o_data_a = 16'b1111110111101000;
            14'h1c38: o_data_a = 16'b1110110010100000;
            14'h1c39: o_data_a = 16'b1110001100001000;
            14'h1c3a: o_data_a = 16'b0000000000000000;
            14'h1c3b: o_data_a = 16'b1111110111001000;
            14'h1c3c: o_data_a = 16'b1111110010100000;
            14'h1c3d: o_data_a = 16'b1110111111001000;
            14'h1c3e: o_data_a = 16'b0000000000000000;
            14'h1c3f: o_data_a = 16'b1111110010101000;
            14'h1c40: o_data_a = 16'b1111110000010000;
            14'h1c41: o_data_a = 16'b1110110010100000;
            14'h1c42: o_data_a = 16'b1111000010001000;
            14'h1c43: o_data_a = 16'b0000000000000000;
            14'h1c44: o_data_a = 16'b1111110010101000;
            14'h1c45: o_data_a = 16'b1111110000010000;
            14'h1c46: o_data_a = 16'b0000000000000001;
            14'h1c47: o_data_a = 16'b1111110111100000;
            14'h1c48: o_data_a = 16'b1110110111100000;
            14'h1c49: o_data_a = 16'b1110110111100000;
            14'h1c4a: o_data_a = 16'b1110001100001000;
            14'h1c4b: o_data_a = 16'b0001101101110101;
            14'h1c4c: o_data_a = 16'b1110101010000111;
            14'h1c4d: o_data_a = 16'b0000000000000001;
            14'h1c4e: o_data_a = 16'b1111110000010000;
            14'h1c4f: o_data_a = 16'b0000000000000100;
            14'h1c50: o_data_a = 16'b1110000010100000;
            14'h1c51: o_data_a = 16'b1111110000010000;
            14'h1c52: o_data_a = 16'b0000000000000000;
            14'h1c53: o_data_a = 16'b1111110111101000;
            14'h1c54: o_data_a = 16'b1110110010100000;
            14'h1c55: o_data_a = 16'b1110001100001000;
            14'h1c56: o_data_a = 16'b0000000000000000;
            14'h1c57: o_data_a = 16'b1111110010101000;
            14'h1c58: o_data_a = 16'b1111110000010000;
            14'h1c59: o_data_a = 16'b0001110001011101;
            14'h1c5a: o_data_a = 16'b1110001100000101;
            14'h1c5b: o_data_a = 16'b0001110001101110;
            14'h1c5c: o_data_a = 16'b1110101010000111;
            14'h1c5d: o_data_a = 16'b0000000000000001;
            14'h1c5e: o_data_a = 16'b1111110000100000;
            14'h1c5f: o_data_a = 16'b1111110000010000;
            14'h1c60: o_data_a = 16'b0000000000000000;
            14'h1c61: o_data_a = 16'b1111110111101000;
            14'h1c62: o_data_a = 16'b1110110010100000;
            14'h1c63: o_data_a = 16'b1110001100001000;
            14'h1c64: o_data_a = 16'b0000000000000000;
            14'h1c65: o_data_a = 16'b1111110010100000;
            14'h1c66: o_data_a = 16'b1111110001010000;
            14'h1c67: o_data_a = 16'b1110011111001000;
            14'h1c68: o_data_a = 16'b0000000000000000;
            14'h1c69: o_data_a = 16'b1111110010101000;
            14'h1c6a: o_data_a = 16'b1111110000010000;
            14'h1c6b: o_data_a = 16'b0000000000000001;
            14'h1c6c: o_data_a = 16'b1111110000100000;
            14'h1c6d: o_data_a = 16'b1110001100001000;
            14'h1c6e: o_data_a = 16'b0000000000000001;
            14'h1c6f: o_data_a = 16'b1111110000100000;
            14'h1c70: o_data_a = 16'b1111110000010000;
            14'h1c71: o_data_a = 16'b0000000000000000;
            14'h1c72: o_data_a = 16'b1111110111101000;
            14'h1c73: o_data_a = 16'b1110110010100000;
            14'h1c74: o_data_a = 16'b1110001100001000;
            14'h1c75: o_data_a = 16'b0000000000110110;
            14'h1c76: o_data_a = 16'b1110101010000111;
            14'h1c77: o_data_a = 16'b0000000000000100;
            14'h1c78: o_data_a = 16'b1110110000010000;
            14'h1c79: o_data_a = 16'b1110001110010000;
            14'h1c7a: o_data_a = 16'b0000000000000000;
            14'h1c7b: o_data_a = 16'b1111110111101000;
            14'h1c7c: o_data_a = 16'b1110110010100000;
            14'h1c7d: o_data_a = 16'b1110101010001000;
            14'h1c7e: o_data_a = 16'b0001110001111001;
            14'h1c7f: o_data_a = 16'b1110001100000001;
            14'h1c80: o_data_a = 16'b0000000000000010;
            14'h1c81: o_data_a = 16'b1111110111100000;
            14'h1c82: o_data_a = 16'b1111110000010000;
            14'h1c83: o_data_a = 16'b0000000000000000;
            14'h1c84: o_data_a = 16'b1111110111101000;
            14'h1c85: o_data_a = 16'b1110110010100000;
            14'h1c86: o_data_a = 16'b1110001100001000;
            14'h1c87: o_data_a = 16'b0000000000000000;
            14'h1c88: o_data_a = 16'b1111110111001000;
            14'h1c89: o_data_a = 16'b1111110010100000;
            14'h1c8a: o_data_a = 16'b1110101010001000;
            14'h1c8b: o_data_a = 16'b0001110010001111;
            14'h1c8c: o_data_a = 16'b1110110000010000;
            14'h1c8d: o_data_a = 16'b0000000000000110;
            14'h1c8e: o_data_a = 16'b1110101010000111;
            14'h1c8f: o_data_a = 16'b0000000000000000;
            14'h1c90: o_data_a = 16'b1111110010101000;
            14'h1c91: o_data_a = 16'b1111110000010000;
            14'h1c92: o_data_a = 16'b0001110010010110;
            14'h1c93: o_data_a = 16'b1110001100000101;
            14'h1c94: o_data_a = 16'b0001110010101101;
            14'h1c95: o_data_a = 16'b1110101010000111;
            14'h1c96: o_data_a = 16'b0000000000000011;
            14'h1c97: o_data_a = 16'b1110110000010000;
            14'h1c98: o_data_a = 16'b0000000000000000;
            14'h1c99: o_data_a = 16'b1111110111101000;
            14'h1c9a: o_data_a = 16'b1110110010100000;
            14'h1c9b: o_data_a = 16'b1110001100001000;
            14'h1c9c: o_data_a = 16'b0000000000000001;
            14'h1c9d: o_data_a = 16'b1110110000010000;
            14'h1c9e: o_data_a = 16'b0000000000001101;
            14'h1c9f: o_data_a = 16'b1110001100001000;
            14'h1ca0: o_data_a = 16'b0110101011011001;
            14'h1ca1: o_data_a = 16'b1110110000010000;
            14'h1ca2: o_data_a = 16'b0000000000001110;
            14'h1ca3: o_data_a = 16'b1110001100001000;
            14'h1ca4: o_data_a = 16'b0001110010101000;
            14'h1ca5: o_data_a = 16'b1110110000010000;
            14'h1ca6: o_data_a = 16'b0000000001011111;
            14'h1ca7: o_data_a = 16'b1110101010000111;
            14'h1ca8: o_data_a = 16'b0000000000000000;
            14'h1ca9: o_data_a = 16'b1111110010101000;
            14'h1caa: o_data_a = 16'b1111110000010000;
            14'h1cab: o_data_a = 16'b0000000000000101;
            14'h1cac: o_data_a = 16'b1110001100001000;
            14'h1cad: o_data_a = 16'b0000000000000010;
            14'h1cae: o_data_a = 16'b1111110000100000;
            14'h1caf: o_data_a = 16'b1111110000010000;
            14'h1cb0: o_data_a = 16'b0000000000000000;
            14'h1cb1: o_data_a = 16'b1111110111101000;
            14'h1cb2: o_data_a = 16'b1110110010100000;
            14'h1cb3: o_data_a = 16'b1110001100001000;
            14'h1cb4: o_data_a = 16'b0000000000000000;
            14'h1cb5: o_data_a = 16'b1111110111001000;
            14'h1cb6: o_data_a = 16'b1111110010100000;
            14'h1cb7: o_data_a = 16'b1110101010001000;
            14'h1cb8: o_data_a = 16'b0001110010111100;
            14'h1cb9: o_data_a = 16'b1110110000010000;
            14'h1cba: o_data_a = 16'b0000000000100110;
            14'h1cbb: o_data_a = 16'b1110101010000111;
            14'h1cbc: o_data_a = 16'b0000000000000010;
            14'h1cbd: o_data_a = 16'b1111110111100000;
            14'h1cbe: o_data_a = 16'b1111110000010000;
            14'h1cbf: o_data_a = 16'b0000000000000000;
            14'h1cc0: o_data_a = 16'b1111110111101000;
            14'h1cc1: o_data_a = 16'b1110110010100000;
            14'h1cc2: o_data_a = 16'b1110001100001000;
            14'h1cc3: o_data_a = 16'b0000000000000000;
            14'h1cc4: o_data_a = 16'b1111110111001000;
            14'h1cc5: o_data_a = 16'b1111110010100000;
            14'h1cc6: o_data_a = 16'b1110101010001000;
            14'h1cc7: o_data_a = 16'b0001110011001011;
            14'h1cc8: o_data_a = 16'b1110110000010000;
            14'h1cc9: o_data_a = 16'b0000000000010110;
            14'h1cca: o_data_a = 16'b1110101010000111;
            14'h1ccb: o_data_a = 16'b0000000000000000;
            14'h1ccc: o_data_a = 16'b1111110010101000;
            14'h1ccd: o_data_a = 16'b1111110000010000;
            14'h1cce: o_data_a = 16'b1110110010100000;
            14'h1ccf: o_data_a = 16'b1111000000001000;
            14'h1cd0: o_data_a = 16'b0000000000000010;
            14'h1cd1: o_data_a = 16'b1111110000100000;
            14'h1cd2: o_data_a = 16'b1111110000010000;
            14'h1cd3: o_data_a = 16'b0000000000000000;
            14'h1cd4: o_data_a = 16'b1111110111101000;
            14'h1cd5: o_data_a = 16'b1110110010100000;
            14'h1cd6: o_data_a = 16'b1110001100001000;
            14'h1cd7: o_data_a = 16'b0000000000000000;
            14'h1cd8: o_data_a = 16'b1111110111001000;
            14'h1cd9: o_data_a = 16'b1111110010100000;
            14'h1cda: o_data_a = 16'b1110101010001000;
            14'h1cdb: o_data_a = 16'b0001110011011111;
            14'h1cdc: o_data_a = 16'b1110110000010000;
            14'h1cdd: o_data_a = 16'b0000000000010110;
            14'h1cde: o_data_a = 16'b1110101010000111;
            14'h1cdf: o_data_a = 16'b0000000000000010;
            14'h1ce0: o_data_a = 16'b1111110111100000;
            14'h1ce1: o_data_a = 16'b1111110000010000;
            14'h1ce2: o_data_a = 16'b0000000000000000;
            14'h1ce3: o_data_a = 16'b1111110111101000;
            14'h1ce4: o_data_a = 16'b1110110010100000;
            14'h1ce5: o_data_a = 16'b1110001100001000;
            14'h1ce6: o_data_a = 16'b0000000000000000;
            14'h1ce7: o_data_a = 16'b1111110111001000;
            14'h1ce8: o_data_a = 16'b1111110010100000;
            14'h1ce9: o_data_a = 16'b1110101010001000;
            14'h1cea: o_data_a = 16'b0001110011101110;
            14'h1ceb: o_data_a = 16'b1110110000010000;
            14'h1cec: o_data_a = 16'b0000000000100110;
            14'h1ced: o_data_a = 16'b1110101010000111;
            14'h1cee: o_data_a = 16'b0000000000000000;
            14'h1cef: o_data_a = 16'b1111110010101000;
            14'h1cf0: o_data_a = 16'b1111110000010000;
            14'h1cf1: o_data_a = 16'b1110110010100000;
            14'h1cf2: o_data_a = 16'b1111000000001000;
            14'h1cf3: o_data_a = 16'b0000000000000000;
            14'h1cf4: o_data_a = 16'b1111110010101000;
            14'h1cf5: o_data_a = 16'b1111110000010000;
            14'h1cf6: o_data_a = 16'b1110110010100000;
            14'h1cf7: o_data_a = 16'b1111010101001000;
            14'h1cf8: o_data_a = 16'b0000000000000000;
            14'h1cf9: o_data_a = 16'b1111110010101000;
            14'h1cfa: o_data_a = 16'b1111110000010000;
            14'h1cfb: o_data_a = 16'b0000000000000001;
            14'h1cfc: o_data_a = 16'b1111110111100000;
            14'h1cfd: o_data_a = 16'b1110110111100000;
            14'h1cfe: o_data_a = 16'b1110001100001000;
            14'h1cff: o_data_a = 16'b0000000000000000;
            14'h1d00: o_data_a = 16'b1111110111001000;
            14'h1d01: o_data_a = 16'b1111110010100000;
            14'h1d02: o_data_a = 16'b1110101010001000;
            14'h1d03: o_data_a = 16'b0000000000010001;
            14'h1d04: o_data_a = 16'b1111110000010000;
            14'h1d05: o_data_a = 16'b0000000000000000;
            14'h1d06: o_data_a = 16'b1111110111101000;
            14'h1d07: o_data_a = 16'b1110110010100000;
            14'h1d08: o_data_a = 16'b1110001100001000;
            14'h1d09: o_data_a = 16'b0000000000000000;
            14'h1d0a: o_data_a = 16'b1111110010101000;
            14'h1d0b: o_data_a = 16'b1111110000010000;
            14'h1d0c: o_data_a = 16'b1110110010100000;
            14'h1d0d: o_data_a = 16'b1111000010001000;
            14'h1d0e: o_data_a = 16'b0000000000000010;
            14'h1d0f: o_data_a = 16'b1111110111100000;
            14'h1d10: o_data_a = 16'b1111110000010000;
            14'h1d11: o_data_a = 16'b0000000000000000;
            14'h1d12: o_data_a = 16'b1111110111101000;
            14'h1d13: o_data_a = 16'b1110110010100000;
            14'h1d14: o_data_a = 16'b1110001100001000;
            14'h1d15: o_data_a = 16'b0000000000000001;
            14'h1d16: o_data_a = 16'b1110110000010000;
            14'h1d17: o_data_a = 16'b0000000000001101;
            14'h1d18: o_data_a = 16'b1110001100001000;
            14'h1d19: o_data_a = 16'b0001101001110110;
            14'h1d1a: o_data_a = 16'b1110110000010000;
            14'h1d1b: o_data_a = 16'b0000000000001110;
            14'h1d1c: o_data_a = 16'b1110001100001000;
            14'h1d1d: o_data_a = 16'b0001110100100001;
            14'h1d1e: o_data_a = 16'b1110110000010000;
            14'h1d1f: o_data_a = 16'b0000000001011111;
            14'h1d20: o_data_a = 16'b1110101010000111;
            14'h1d21: o_data_a = 16'b0000000000000000;
            14'h1d22: o_data_a = 16'b1111110010101000;
            14'h1d23: o_data_a = 16'b1111110000010000;
            14'h1d24: o_data_a = 16'b0000000000000101;
            14'h1d25: o_data_a = 16'b1110001100001000;
            14'h1d26: o_data_a = 16'b0000000000000000;
            14'h1d27: o_data_a = 16'b1111110010101000;
            14'h1d28: o_data_a = 16'b1111110000010000;
            14'h1d29: o_data_a = 16'b0000000000000100;
            14'h1d2a: o_data_a = 16'b1110001100001000;
            14'h1d2b: o_data_a = 16'b0000000000000101;
            14'h1d2c: o_data_a = 16'b1111110000010000;
            14'h1d2d: o_data_a = 16'b0000000000000000;
            14'h1d2e: o_data_a = 16'b1111110111101000;
            14'h1d2f: o_data_a = 16'b1110110010100000;
            14'h1d30: o_data_a = 16'b1110001100001000;
            14'h1d31: o_data_a = 16'b0000000000000000;
            14'h1d32: o_data_a = 16'b1111110010101000;
            14'h1d33: o_data_a = 16'b1111110000010000;
            14'h1d34: o_data_a = 16'b0000000000000100;
            14'h1d35: o_data_a = 16'b1111110000100000;
            14'h1d36: o_data_a = 16'b1110001100001000;
            14'h1d37: o_data_a = 16'b0000000000000010;
            14'h1d38: o_data_a = 16'b1111110000100000;
            14'h1d39: o_data_a = 16'b1111110000010000;
            14'h1d3a: o_data_a = 16'b0000000000000000;
            14'h1d3b: o_data_a = 16'b1111110111101000;
            14'h1d3c: o_data_a = 16'b1110110010100000;
            14'h1d3d: o_data_a = 16'b1110001100001000;
            14'h1d3e: o_data_a = 16'b0000000000000001;
            14'h1d3f: o_data_a = 16'b1110110000010000;
            14'h1d40: o_data_a = 16'b0000000000001101;
            14'h1d41: o_data_a = 16'b1110001100001000;
            14'h1d42: o_data_a = 16'b0001101001110110;
            14'h1d43: o_data_a = 16'b1110110000010000;
            14'h1d44: o_data_a = 16'b0000000000001110;
            14'h1d45: o_data_a = 16'b1110001100001000;
            14'h1d46: o_data_a = 16'b0001110101001010;
            14'h1d47: o_data_a = 16'b1110110000010000;
            14'h1d48: o_data_a = 16'b0000000001011111;
            14'h1d49: o_data_a = 16'b1110101010000111;
            14'h1d4a: o_data_a = 16'b0000000000000000;
            14'h1d4b: o_data_a = 16'b1111110010101000;
            14'h1d4c: o_data_a = 16'b1111110000010000;
            14'h1d4d: o_data_a = 16'b0000000000000010;
            14'h1d4e: o_data_a = 16'b1111110000100000;
            14'h1d4f: o_data_a = 16'b1110001100001000;
            14'h1d50: o_data_a = 16'b0000000000000001;
            14'h1d51: o_data_a = 16'b1111110000010000;
            14'h1d52: o_data_a = 16'b0000000000000011;
            14'h1d53: o_data_a = 16'b1110000010100000;
            14'h1d54: o_data_a = 16'b1111110000010000;
            14'h1d55: o_data_a = 16'b0000000000000000;
            14'h1d56: o_data_a = 16'b1111110111101000;
            14'h1d57: o_data_a = 16'b1110110010100000;
            14'h1d58: o_data_a = 16'b1110001100001000;
            14'h1d59: o_data_a = 16'b0000000000000000;
            14'h1d5a: o_data_a = 16'b1111110010100000;
            14'h1d5b: o_data_a = 16'b1111110001001000;
            14'h1d5c: o_data_a = 16'b0000000000000000;
            14'h1d5d: o_data_a = 16'b1111110010100000;
            14'h1d5e: o_data_a = 16'b1111110001001000;
            14'h1d5f: o_data_a = 16'b0000000000000000;
            14'h1d60: o_data_a = 16'b1111110010101000;
            14'h1d61: o_data_a = 16'b1111110000010000;
            14'h1d62: o_data_a = 16'b0001111010100001;
            14'h1d63: o_data_a = 16'b1110001100000101;
            14'h1d64: o_data_a = 16'b0111111111111111;
            14'h1d65: o_data_a = 16'b1110110000010000;
            14'h1d66: o_data_a = 16'b0000000000000000;
            14'h1d67: o_data_a = 16'b1111110111101000;
            14'h1d68: o_data_a = 16'b1110110010100000;
            14'h1d69: o_data_a = 16'b1110001100001000;
            14'h1d6a: o_data_a = 16'b0000000000000001;
            14'h1d6b: o_data_a = 16'b1111110000100000;
            14'h1d6c: o_data_a = 16'b1111110000010000;
            14'h1d6d: o_data_a = 16'b0000000000000000;
            14'h1d6e: o_data_a = 16'b1111110111101000;
            14'h1d6f: o_data_a = 16'b1110110010100000;
            14'h1d70: o_data_a = 16'b1110001100001000;
            14'h1d71: o_data_a = 16'b0000000000010001;
            14'h1d72: o_data_a = 16'b1111110000010000;
            14'h1d73: o_data_a = 16'b0000000000000000;
            14'h1d74: o_data_a = 16'b1111110111101000;
            14'h1d75: o_data_a = 16'b1110110010100000;
            14'h1d76: o_data_a = 16'b1110001100001000;
            14'h1d77: o_data_a = 16'b0000000000000000;
            14'h1d78: o_data_a = 16'b1111110010101000;
            14'h1d79: o_data_a = 16'b1111110000010000;
            14'h1d7a: o_data_a = 16'b1110110010100000;
            14'h1d7b: o_data_a = 16'b1111000010001000;
            14'h1d7c: o_data_a = 16'b0000000000000000;
            14'h1d7d: o_data_a = 16'b1111110010101000;
            14'h1d7e: o_data_a = 16'b1111110000010000;
            14'h1d7f: o_data_a = 16'b0000000000000100;
            14'h1d80: o_data_a = 16'b1110001100001000;
            14'h1d81: o_data_a = 16'b0000000000000100;
            14'h1d82: o_data_a = 16'b1111110000100000;
            14'h1d83: o_data_a = 16'b1111110000010000;
            14'h1d84: o_data_a = 16'b0000000000000000;
            14'h1d85: o_data_a = 16'b1111110111101000;
            14'h1d86: o_data_a = 16'b1110110010100000;
            14'h1d87: o_data_a = 16'b1110001100001000;
            14'h1d88: o_data_a = 16'b0000000000000000;
            14'h1d89: o_data_a = 16'b1111110010101000;
            14'h1d8a: o_data_a = 16'b1111110000010000;
            14'h1d8b: o_data_a = 16'b1110110010100000;
            14'h1d8c: o_data_a = 16'b1111000111001000;
            14'h1d8d: o_data_a = 16'b0000000000000001;
            14'h1d8e: o_data_a = 16'b1111110000100000;
            14'h1d8f: o_data_a = 16'b1111110000010000;
            14'h1d90: o_data_a = 16'b0000000000000000;
            14'h1d91: o_data_a = 16'b1111110111101000;
            14'h1d92: o_data_a = 16'b1110110010100000;
            14'h1d93: o_data_a = 16'b1110001100001000;
            14'h1d94: o_data_a = 16'b0000000000010001;
            14'h1d95: o_data_a = 16'b1111110000010000;
            14'h1d96: o_data_a = 16'b0000000000000000;
            14'h1d97: o_data_a = 16'b1111110111101000;
            14'h1d98: o_data_a = 16'b1110110010100000;
            14'h1d99: o_data_a = 16'b1110001100001000;
            14'h1d9a: o_data_a = 16'b0000000000000000;
            14'h1d9b: o_data_a = 16'b1111110010101000;
            14'h1d9c: o_data_a = 16'b1111110000010000;
            14'h1d9d: o_data_a = 16'b1110110010100000;
            14'h1d9e: o_data_a = 16'b1111000010001000;
            14'h1d9f: o_data_a = 16'b0000000000000000;
            14'h1da0: o_data_a = 16'b1111110010101000;
            14'h1da1: o_data_a = 16'b1111110000010000;
            14'h1da2: o_data_a = 16'b0000000000000100;
            14'h1da3: o_data_a = 16'b1110001100001000;
            14'h1da4: o_data_a = 16'b0000000000000100;
            14'h1da5: o_data_a = 16'b1111110000100000;
            14'h1da6: o_data_a = 16'b1111110000010000;
            14'h1da7: o_data_a = 16'b0000000000000000;
            14'h1da8: o_data_a = 16'b1111110111101000;
            14'h1da9: o_data_a = 16'b1110110010100000;
            14'h1daa: o_data_a = 16'b1110001100001000;
            14'h1dab: o_data_a = 16'b0001110110101111;
            14'h1dac: o_data_a = 16'b1110110000010000;
            14'h1dad: o_data_a = 16'b0000000000100110;
            14'h1dae: o_data_a = 16'b1110101010000111;
            14'h1daf: o_data_a = 16'b0000000000000000;
            14'h1db0: o_data_a = 16'b1111110010101000;
            14'h1db1: o_data_a = 16'b1111110000010000;
            14'h1db2: o_data_a = 16'b0000000000000001;
            14'h1db3: o_data_a = 16'b1111110111100000;
            14'h1db4: o_data_a = 16'b1110110111100000;
            14'h1db5: o_data_a = 16'b1110110111100000;
            14'h1db6: o_data_a = 16'b1110001100001000;
            14'h1db7: o_data_a = 16'b0000000000000001;
            14'h1db8: o_data_a = 16'b1111110000010000;
            14'h1db9: o_data_a = 16'b0000000000000011;
            14'h1dba: o_data_a = 16'b1110000010100000;
            14'h1dbb: o_data_a = 16'b1111110000010000;
            14'h1dbc: o_data_a = 16'b0000000000000000;
            14'h1dbd: o_data_a = 16'b1111110111101000;
            14'h1dbe: o_data_a = 16'b1110110010100000;
            14'h1dbf: o_data_a = 16'b1110001100001000;
            14'h1dc0: o_data_a = 16'b0000000000000000;
            14'h1dc1: o_data_a = 16'b1111110010100000;
            14'h1dc2: o_data_a = 16'b1111110001001000;
            14'h1dc3: o_data_a = 16'b0000000000000000;
            14'h1dc4: o_data_a = 16'b1111110010101000;
            14'h1dc5: o_data_a = 16'b1111110000010000;
            14'h1dc6: o_data_a = 16'b0001110111001010;
            14'h1dc7: o_data_a = 16'b1110001100000101;
            14'h1dc8: o_data_a = 16'b0001111010011111;
            14'h1dc9: o_data_a = 16'b1110101010000111;
            14'h1dca: o_data_a = 16'b0000000000000001;
            14'h1dcb: o_data_a = 16'b1111110000100000;
            14'h1dcc: o_data_a = 16'b1111110000010000;
            14'h1dcd: o_data_a = 16'b0000000000000000;
            14'h1dce: o_data_a = 16'b1111110111101000;
            14'h1dcf: o_data_a = 16'b1110110010100000;
            14'h1dd0: o_data_a = 16'b1110001100001000;
            14'h1dd1: o_data_a = 16'b0000000000000000;
            14'h1dd2: o_data_a = 16'b1111110111001000;
            14'h1dd3: o_data_a = 16'b1111110010100000;
            14'h1dd4: o_data_a = 16'b1110111111001000;
            14'h1dd5: o_data_a = 16'b0000000000000000;
            14'h1dd6: o_data_a = 16'b1111110010101000;
            14'h1dd7: o_data_a = 16'b1111110000010000;
            14'h1dd8: o_data_a = 16'b1110110010100000;
            14'h1dd9: o_data_a = 16'b1111000010001000;
            14'h1dda: o_data_a = 16'b0000000000010001;
            14'h1ddb: o_data_a = 16'b1111110000010000;
            14'h1ddc: o_data_a = 16'b0000000000000000;
            14'h1ddd: o_data_a = 16'b1111110111101000;
            14'h1dde: o_data_a = 16'b1110110010100000;
            14'h1ddf: o_data_a = 16'b1110001100001000;
            14'h1de0: o_data_a = 16'b0000000000000000;
            14'h1de1: o_data_a = 16'b1111110010101000;
            14'h1de2: o_data_a = 16'b1111110000010000;
            14'h1de3: o_data_a = 16'b1110110010100000;
            14'h1de4: o_data_a = 16'b1111000010001000;
            14'h1de5: o_data_a = 16'b0000000000000001;
            14'h1de6: o_data_a = 16'b1111110000100000;
            14'h1de7: o_data_a = 16'b1111110000010000;
            14'h1de8: o_data_a = 16'b0000000000000000;
            14'h1de9: o_data_a = 16'b1111110111101000;
            14'h1dea: o_data_a = 16'b1110110010100000;
            14'h1deb: o_data_a = 16'b1110001100001000;
            14'h1dec: o_data_a = 16'b0000000000010001;
            14'h1ded: o_data_a = 16'b1111110000010000;
            14'h1dee: o_data_a = 16'b0000000000000000;
            14'h1def: o_data_a = 16'b1111110111101000;
            14'h1df0: o_data_a = 16'b1110110010100000;
            14'h1df1: o_data_a = 16'b1110001100001000;
            14'h1df2: o_data_a = 16'b0000000000000000;
            14'h1df3: o_data_a = 16'b1111110010101000;
            14'h1df4: o_data_a = 16'b1111110000010000;
            14'h1df5: o_data_a = 16'b1110110010100000;
            14'h1df6: o_data_a = 16'b1111000010001000;
            14'h1df7: o_data_a = 16'b0000000000000000;
            14'h1df8: o_data_a = 16'b1111110010101000;
            14'h1df9: o_data_a = 16'b1111110000010000;
            14'h1dfa: o_data_a = 16'b0000000000000100;
            14'h1dfb: o_data_a = 16'b1110001100001000;
            14'h1dfc: o_data_a = 16'b0000000000000100;
            14'h1dfd: o_data_a = 16'b1111110000100000;
            14'h1dfe: o_data_a = 16'b1111110000010000;
            14'h1dff: o_data_a = 16'b0000000000000000;
            14'h1e00: o_data_a = 16'b1111110111101000;
            14'h1e01: o_data_a = 16'b1110110010100000;
            14'h1e02: o_data_a = 16'b1110001100001000;
            14'h1e03: o_data_a = 16'b0000000000000001;
            14'h1e04: o_data_a = 16'b1111110000100000;
            14'h1e05: o_data_a = 16'b1111110000010000;
            14'h1e06: o_data_a = 16'b0000000000000000;
            14'h1e07: o_data_a = 16'b1111110111101000;
            14'h1e08: o_data_a = 16'b1110110010100000;
            14'h1e09: o_data_a = 16'b1110001100001000;
            14'h1e0a: o_data_a = 16'b0000000000010001;
            14'h1e0b: o_data_a = 16'b1111110000010000;
            14'h1e0c: o_data_a = 16'b0000000000000000;
            14'h1e0d: o_data_a = 16'b1111110111101000;
            14'h1e0e: o_data_a = 16'b1110110010100000;
            14'h1e0f: o_data_a = 16'b1110001100001000;
            14'h1e10: o_data_a = 16'b0000000000000000;
            14'h1e11: o_data_a = 16'b1111110010101000;
            14'h1e12: o_data_a = 16'b1111110000010000;
            14'h1e13: o_data_a = 16'b1110110010100000;
            14'h1e14: o_data_a = 16'b1111000010001000;
            14'h1e15: o_data_a = 16'b0000000000000000;
            14'h1e16: o_data_a = 16'b1111110010101000;
            14'h1e17: o_data_a = 16'b1111110000010000;
            14'h1e18: o_data_a = 16'b0000000000000100;
            14'h1e19: o_data_a = 16'b1110001100001000;
            14'h1e1a: o_data_a = 16'b0000000000000100;
            14'h1e1b: o_data_a = 16'b1111110000100000;
            14'h1e1c: o_data_a = 16'b1111110000010000;
            14'h1e1d: o_data_a = 16'b0000000000000000;
            14'h1e1e: o_data_a = 16'b1111110111101000;
            14'h1e1f: o_data_a = 16'b1110110010100000;
            14'h1e20: o_data_a = 16'b1110001100001000;
            14'h1e21: o_data_a = 16'b0000000000000000;
            14'h1e22: o_data_a = 16'b1111110010101000;
            14'h1e23: o_data_a = 16'b1111110000010000;
            14'h1e24: o_data_a = 16'b1110110010100000;
            14'h1e25: o_data_a = 16'b1111000010001000;
            14'h1e26: o_data_a = 16'b0000000000000000;
            14'h1e27: o_data_a = 16'b1111110010101000;
            14'h1e28: o_data_a = 16'b1111110000010000;
            14'h1e29: o_data_a = 16'b0000000000000101;
            14'h1e2a: o_data_a = 16'b1110001100001000;
            14'h1e2b: o_data_a = 16'b0000000000000000;
            14'h1e2c: o_data_a = 16'b1111110010101000;
            14'h1e2d: o_data_a = 16'b1111110000010000;
            14'h1e2e: o_data_a = 16'b0000000000000100;
            14'h1e2f: o_data_a = 16'b1110001100001000;
            14'h1e30: o_data_a = 16'b0000000000000101;
            14'h1e31: o_data_a = 16'b1111110000010000;
            14'h1e32: o_data_a = 16'b0000000000000000;
            14'h1e33: o_data_a = 16'b1111110111101000;
            14'h1e34: o_data_a = 16'b1110110010100000;
            14'h1e35: o_data_a = 16'b1110001100001000;
            14'h1e36: o_data_a = 16'b0000000000000000;
            14'h1e37: o_data_a = 16'b1111110010101000;
            14'h1e38: o_data_a = 16'b1111110000010000;
            14'h1e39: o_data_a = 16'b0000000000000100;
            14'h1e3a: o_data_a = 16'b1111110000100000;
            14'h1e3b: o_data_a = 16'b1110001100001000;
            14'h1e3c: o_data_a = 16'b0000000000000001;
            14'h1e3d: o_data_a = 16'b1111110000100000;
            14'h1e3e: o_data_a = 16'b1111110000010000;
            14'h1e3f: o_data_a = 16'b0000000000000000;
            14'h1e40: o_data_a = 16'b1111110111101000;
            14'h1e41: o_data_a = 16'b1110110010100000;
            14'h1e42: o_data_a = 16'b1110001100001000;
            14'h1e43: o_data_a = 16'b0000000000000000;
            14'h1e44: o_data_a = 16'b1111110111001000;
            14'h1e45: o_data_a = 16'b1111110010100000;
            14'h1e46: o_data_a = 16'b1110111111001000;
            14'h1e47: o_data_a = 16'b0000000000000000;
            14'h1e48: o_data_a = 16'b1111110010101000;
            14'h1e49: o_data_a = 16'b1111110000010000;
            14'h1e4a: o_data_a = 16'b1110110010100000;
            14'h1e4b: o_data_a = 16'b1111000010001000;
            14'h1e4c: o_data_a = 16'b0000000000010001;
            14'h1e4d: o_data_a = 16'b1111110000010000;
            14'h1e4e: o_data_a = 16'b0000000000000000;
            14'h1e4f: o_data_a = 16'b1111110111101000;
            14'h1e50: o_data_a = 16'b1110110010100000;
            14'h1e51: o_data_a = 16'b1110001100001000;
            14'h1e52: o_data_a = 16'b0000000000000000;
            14'h1e53: o_data_a = 16'b1111110010101000;
            14'h1e54: o_data_a = 16'b1111110000010000;
            14'h1e55: o_data_a = 16'b1110110010100000;
            14'h1e56: o_data_a = 16'b1111000010001000;
            14'h1e57: o_data_a = 16'b0000000000000000;
            14'h1e58: o_data_a = 16'b1111110010101000;
            14'h1e59: o_data_a = 16'b1111110000010000;
            14'h1e5a: o_data_a = 16'b0000000000000100;
            14'h1e5b: o_data_a = 16'b1110001100001000;
            14'h1e5c: o_data_a = 16'b0000000000000100;
            14'h1e5d: o_data_a = 16'b1111110000100000;
            14'h1e5e: o_data_a = 16'b1111110000010000;
            14'h1e5f: o_data_a = 16'b0000000000000000;
            14'h1e60: o_data_a = 16'b1111110111101000;
            14'h1e61: o_data_a = 16'b1110110010100000;
            14'h1e62: o_data_a = 16'b1110001100001000;
            14'h1e63: o_data_a = 16'b0000000000000010;
            14'h1e64: o_data_a = 16'b1111110000100000;
            14'h1e65: o_data_a = 16'b1111110000010000;
            14'h1e66: o_data_a = 16'b0000000000000000;
            14'h1e67: o_data_a = 16'b1111110111101000;
            14'h1e68: o_data_a = 16'b1110110010100000;
            14'h1e69: o_data_a = 16'b1110001100001000;
            14'h1e6a: o_data_a = 16'b0001111001101110;
            14'h1e6b: o_data_a = 16'b1110110000010000;
            14'h1e6c: o_data_a = 16'b0000000000010110;
            14'h1e6d: o_data_a = 16'b1110101010000111;
            14'h1e6e: o_data_a = 16'b0000000000000000;
            14'h1e6f: o_data_a = 16'b1111110010101000;
            14'h1e70: o_data_a = 16'b1111110000010000;
            14'h1e71: o_data_a = 16'b0000000000000001;
            14'h1e72: o_data_a = 16'b1111110111100000;
            14'h1e73: o_data_a = 16'b1110110111100000;
            14'h1e74: o_data_a = 16'b1110110111100000;
            14'h1e75: o_data_a = 16'b1110001100001000;
            14'h1e76: o_data_a = 16'b0000000000000001;
            14'h1e77: o_data_a = 16'b1111110000010000;
            14'h1e78: o_data_a = 16'b0000000000000011;
            14'h1e79: o_data_a = 16'b1110000010100000;
            14'h1e7a: o_data_a = 16'b1111110000010000;
            14'h1e7b: o_data_a = 16'b0000000000000000;
            14'h1e7c: o_data_a = 16'b1111110111101000;
            14'h1e7d: o_data_a = 16'b1110110010100000;
            14'h1e7e: o_data_a = 16'b1110001100001000;
            14'h1e7f: o_data_a = 16'b0000000000000000;
            14'h1e80: o_data_a = 16'b1111110010100000;
            14'h1e81: o_data_a = 16'b1111110001001000;
            14'h1e82: o_data_a = 16'b0000000000000000;
            14'h1e83: o_data_a = 16'b1111110010101000;
            14'h1e84: o_data_a = 16'b1111110000010000;
            14'h1e85: o_data_a = 16'b0001111010001001;
            14'h1e86: o_data_a = 16'b1110001100000101;
            14'h1e87: o_data_a = 16'b0001111010011111;
            14'h1e88: o_data_a = 16'b1110101010000111;
            14'h1e89: o_data_a = 16'b0000000000000001;
            14'h1e8a: o_data_a = 16'b1111110000100000;
            14'h1e8b: o_data_a = 16'b1111110000010000;
            14'h1e8c: o_data_a = 16'b0000000000000000;
            14'h1e8d: o_data_a = 16'b1111110111101000;
            14'h1e8e: o_data_a = 16'b1110110010100000;
            14'h1e8f: o_data_a = 16'b1110001100001000;
            14'h1e90: o_data_a = 16'b0000000000000000;
            14'h1e91: o_data_a = 16'b1111110111001000;
            14'h1e92: o_data_a = 16'b1111110010100000;
            14'h1e93: o_data_a = 16'b1110111111001000;
            14'h1e94: o_data_a = 16'b0000000000000000;
            14'h1e95: o_data_a = 16'b1111110010101000;
            14'h1e96: o_data_a = 16'b1111110000010000;
            14'h1e97: o_data_a = 16'b1110110010100000;
            14'h1e98: o_data_a = 16'b1111000010001000;
            14'h1e99: o_data_a = 16'b0000000000000000;
            14'h1e9a: o_data_a = 16'b1111110010101000;
            14'h1e9b: o_data_a = 16'b1111110000010000;
            14'h1e9c: o_data_a = 16'b0000000000000001;
            14'h1e9d: o_data_a = 16'b1111110000100000;
            14'h1e9e: o_data_a = 16'b1110001100001000;
            14'h1e9f: o_data_a = 16'b0001110101010000;
            14'h1ea0: o_data_a = 16'b1110101010000111;
            14'h1ea1: o_data_a = 16'b0000000000000001;
            14'h1ea2: o_data_a = 16'b1111110000100000;
            14'h1ea3: o_data_a = 16'b1111110000010000;
            14'h1ea4: o_data_a = 16'b0000000000000000;
            14'h1ea5: o_data_a = 16'b1111110111101000;
            14'h1ea6: o_data_a = 16'b1110110010100000;
            14'h1ea7: o_data_a = 16'b1110001100001000;
            14'h1ea8: o_data_a = 16'b0000000000000000;
            14'h1ea9: o_data_a = 16'b1111110111001000;
            14'h1eaa: o_data_a = 16'b1111110010100000;
            14'h1eab: o_data_a = 16'b1110111111001000;
            14'h1eac: o_data_a = 16'b0000000000000000;
            14'h1ead: o_data_a = 16'b1111110010100000;
            14'h1eae: o_data_a = 16'b1111110001010000;
            14'h1eaf: o_data_a = 16'b1110011111001000;
            14'h1eb0: o_data_a = 16'b0001111010110100;
            14'h1eb1: o_data_a = 16'b1110110000010000;
            14'h1eb2: o_data_a = 16'b0000000000010110;
            14'h1eb3: o_data_a = 16'b1110101010000111;
            14'h1eb4: o_data_a = 16'b0000000000000000;
            14'h1eb5: o_data_a = 16'b1111110010100000;
            14'h1eb6: o_data_a = 16'b1111110001001000;
            14'h1eb7: o_data_a = 16'b0000000000000000;
            14'h1eb8: o_data_a = 16'b1111110010101000;
            14'h1eb9: o_data_a = 16'b1111110000010000;
            14'h1eba: o_data_a = 16'b0001111101100111;
            14'h1ebb: o_data_a = 16'b1110001100000101;
            14'h1ebc: o_data_a = 16'b0000000000000001;
            14'h1ebd: o_data_a = 16'b1111110000100000;
            14'h1ebe: o_data_a = 16'b1111110000010000;
            14'h1ebf: o_data_a = 16'b0000000000000000;
            14'h1ec0: o_data_a = 16'b1111110111101000;
            14'h1ec1: o_data_a = 16'b1110110010100000;
            14'h1ec2: o_data_a = 16'b1110001100001000;
            14'h1ec3: o_data_a = 16'b0000000000010001;
            14'h1ec4: o_data_a = 16'b1111110000010000;
            14'h1ec5: o_data_a = 16'b0000000000000000;
            14'h1ec6: o_data_a = 16'b1111110111101000;
            14'h1ec7: o_data_a = 16'b1110110010100000;
            14'h1ec8: o_data_a = 16'b1110001100001000;
            14'h1ec9: o_data_a = 16'b0000000000000000;
            14'h1eca: o_data_a = 16'b1111110010101000;
            14'h1ecb: o_data_a = 16'b1111110000010000;
            14'h1ecc: o_data_a = 16'b1110110010100000;
            14'h1ecd: o_data_a = 16'b1111000010001000;
            14'h1ece: o_data_a = 16'b0000000000000000;
            14'h1ecf: o_data_a = 16'b1111110010101000;
            14'h1ed0: o_data_a = 16'b1111110000010000;
            14'h1ed1: o_data_a = 16'b0000000000000100;
            14'h1ed2: o_data_a = 16'b1110001100001000;
            14'h1ed3: o_data_a = 16'b0000000000000100;
            14'h1ed4: o_data_a = 16'b1111110000100000;
            14'h1ed5: o_data_a = 16'b1111110000010000;
            14'h1ed6: o_data_a = 16'b0000000000000000;
            14'h1ed7: o_data_a = 16'b1111110111101000;
            14'h1ed8: o_data_a = 16'b1110110010100000;
            14'h1ed9: o_data_a = 16'b1110001100001000;
            14'h1eda: o_data_a = 16'b0000000000000010;
            14'h1edb: o_data_a = 16'b1111110000100000;
            14'h1edc: o_data_a = 16'b1111110000010000;
            14'h1edd: o_data_a = 16'b0000000000000000;
            14'h1ede: o_data_a = 16'b1111110111101000;
            14'h1edf: o_data_a = 16'b1110110010100000;
            14'h1ee0: o_data_a = 16'b1110001100001000;
            14'h1ee1: o_data_a = 16'b0001111011100101;
            14'h1ee2: o_data_a = 16'b1110110000010000;
            14'h1ee3: o_data_a = 16'b0000000000010110;
            14'h1ee4: o_data_a = 16'b1110101010000111;
            14'h1ee5: o_data_a = 16'b0000000000000000;
            14'h1ee6: o_data_a = 16'b1111110010100000;
            14'h1ee7: o_data_a = 16'b1111110001001000;
            14'h1ee8: o_data_a = 16'b0000000000000000;
            14'h1ee9: o_data_a = 16'b1111110010101000;
            14'h1eea: o_data_a = 16'b1111110000010000;
            14'h1eeb: o_data_a = 16'b0001111011101111;
            14'h1eec: o_data_a = 16'b1110001100000101;
            14'h1eed: o_data_a = 16'b0001111101001111;
            14'h1eee: o_data_a = 16'b1110101010000111;
            14'h1eef: o_data_a = 16'b0000000000000001;
            14'h1ef0: o_data_a = 16'b1111110111100000;
            14'h1ef1: o_data_a = 16'b1111110000010000;
            14'h1ef2: o_data_a = 16'b0000000000000000;
            14'h1ef3: o_data_a = 16'b1111110111101000;
            14'h1ef4: o_data_a = 16'b1110110010100000;
            14'h1ef5: o_data_a = 16'b1110001100001000;
            14'h1ef6: o_data_a = 16'b0000000000000001;
            14'h1ef7: o_data_a = 16'b1111110000100000;
            14'h1ef8: o_data_a = 16'b1111110000010000;
            14'h1ef9: o_data_a = 16'b0000000000000000;
            14'h1efa: o_data_a = 16'b1111110111101000;
            14'h1efb: o_data_a = 16'b1110110010100000;
            14'h1efc: o_data_a = 16'b1110001100001000;
            14'h1efd: o_data_a = 16'b0000000000010010;
            14'h1efe: o_data_a = 16'b1111110000010000;
            14'h1eff: o_data_a = 16'b0000000000000000;
            14'h1f00: o_data_a = 16'b1111110111101000;
            14'h1f01: o_data_a = 16'b1110110010100000;
            14'h1f02: o_data_a = 16'b1110001100001000;
            14'h1f03: o_data_a = 16'b0000000000000000;
            14'h1f04: o_data_a = 16'b1111110010101000;
            14'h1f05: o_data_a = 16'b1111110000010000;
            14'h1f06: o_data_a = 16'b1110110010100000;
            14'h1f07: o_data_a = 16'b1111000010001000;
            14'h1f08: o_data_a = 16'b0000000000000000;
            14'h1f09: o_data_a = 16'b1111110010101000;
            14'h1f0a: o_data_a = 16'b1111110000010000;
            14'h1f0b: o_data_a = 16'b0000000000000100;
            14'h1f0c: o_data_a = 16'b1110001100001000;
            14'h1f0d: o_data_a = 16'b0000000000000100;
            14'h1f0e: o_data_a = 16'b1111110000100000;
            14'h1f0f: o_data_a = 16'b1111110000010000;
            14'h1f10: o_data_a = 16'b0000000000000000;
            14'h1f11: o_data_a = 16'b1111110111101000;
            14'h1f12: o_data_a = 16'b1110110010100000;
            14'h1f13: o_data_a = 16'b1110001100001000;
            14'h1f14: o_data_a = 16'b0000000000000000;
            14'h1f15: o_data_a = 16'b1111110010101000;
            14'h1f16: o_data_a = 16'b1111110000010000;
            14'h1f17: o_data_a = 16'b1110110010100000;
            14'h1f18: o_data_a = 16'b1111000010001000;
            14'h1f19: o_data_a = 16'b0000000000000000;
            14'h1f1a: o_data_a = 16'b1111110010101000;
            14'h1f1b: o_data_a = 16'b1111110000010000;
            14'h1f1c: o_data_a = 16'b0000000000000001;
            14'h1f1d: o_data_a = 16'b1111110111100000;
            14'h1f1e: o_data_a = 16'b1110001100001000;
            14'h1f1f: o_data_a = 16'b0000000000000010;
            14'h1f20: o_data_a = 16'b1111110000100000;
            14'h1f21: o_data_a = 16'b1111110000010000;
            14'h1f22: o_data_a = 16'b0000000000000000;
            14'h1f23: o_data_a = 16'b1111110111101000;
            14'h1f24: o_data_a = 16'b1110110010100000;
            14'h1f25: o_data_a = 16'b1110001100001000;
            14'h1f26: o_data_a = 16'b0000000000000001;
            14'h1f27: o_data_a = 16'b1111110000100000;
            14'h1f28: o_data_a = 16'b1111110000010000;
            14'h1f29: o_data_a = 16'b0000000000000000;
            14'h1f2a: o_data_a = 16'b1111110111101000;
            14'h1f2b: o_data_a = 16'b1110110010100000;
            14'h1f2c: o_data_a = 16'b1110001100001000;
            14'h1f2d: o_data_a = 16'b0000000000010001;
            14'h1f2e: o_data_a = 16'b1111110000010000;
            14'h1f2f: o_data_a = 16'b0000000000000000;
            14'h1f30: o_data_a = 16'b1111110111101000;
            14'h1f31: o_data_a = 16'b1110110010100000;
            14'h1f32: o_data_a = 16'b1110001100001000;
            14'h1f33: o_data_a = 16'b0000000000000000;
            14'h1f34: o_data_a = 16'b1111110010101000;
            14'h1f35: o_data_a = 16'b1111110000010000;
            14'h1f36: o_data_a = 16'b1110110010100000;
            14'h1f37: o_data_a = 16'b1111000010001000;
            14'h1f38: o_data_a = 16'b0000000000000000;
            14'h1f39: o_data_a = 16'b1111110010101000;
            14'h1f3a: o_data_a = 16'b1111110000010000;
            14'h1f3b: o_data_a = 16'b0000000000000100;
            14'h1f3c: o_data_a = 16'b1110001100001000;
            14'h1f3d: o_data_a = 16'b0000000000000100;
            14'h1f3e: o_data_a = 16'b1111110000100000;
            14'h1f3f: o_data_a = 16'b1111110000010000;
            14'h1f40: o_data_a = 16'b0000000000000000;
            14'h1f41: o_data_a = 16'b1111110111101000;
            14'h1f42: o_data_a = 16'b1110110010100000;
            14'h1f43: o_data_a = 16'b1110001100001000;
            14'h1f44: o_data_a = 16'b0000000000000000;
            14'h1f45: o_data_a = 16'b1111110010101000;
            14'h1f46: o_data_a = 16'b1111110000010000;
            14'h1f47: o_data_a = 16'b1110110010100000;
            14'h1f48: o_data_a = 16'b1111000111001000;
            14'h1f49: o_data_a = 16'b0000000000000000;
            14'h1f4a: o_data_a = 16'b1111110010101000;
            14'h1f4b: o_data_a = 16'b1111110000010000;
            14'h1f4c: o_data_a = 16'b0000000000000010;
            14'h1f4d: o_data_a = 16'b1111110000100000;
            14'h1f4e: o_data_a = 16'b1110001100001000;
            14'h1f4f: o_data_a = 16'b0000000000000001;
            14'h1f50: o_data_a = 16'b1111110000100000;
            14'h1f51: o_data_a = 16'b1111110000010000;
            14'h1f52: o_data_a = 16'b0000000000000000;
            14'h1f53: o_data_a = 16'b1111110111101000;
            14'h1f54: o_data_a = 16'b1110110010100000;
            14'h1f55: o_data_a = 16'b1110001100001000;
            14'h1f56: o_data_a = 16'b0000000000000000;
            14'h1f57: o_data_a = 16'b1111110111001000;
            14'h1f58: o_data_a = 16'b1111110010100000;
            14'h1f59: o_data_a = 16'b1110111111001000;
            14'h1f5a: o_data_a = 16'b0000000000000000;
            14'h1f5b: o_data_a = 16'b1111110010101000;
            14'h1f5c: o_data_a = 16'b1111110000010000;
            14'h1f5d: o_data_a = 16'b1110110010100000;
            14'h1f5e: o_data_a = 16'b1111000111001000;
            14'h1f5f: o_data_a = 16'b0000000000000000;
            14'h1f60: o_data_a = 16'b1111110010101000;
            14'h1f61: o_data_a = 16'b1111110000010000;
            14'h1f62: o_data_a = 16'b0000000000000001;
            14'h1f63: o_data_a = 16'b1111110000100000;
            14'h1f64: o_data_a = 16'b1110001100001000;
            14'h1f65: o_data_a = 16'b0001111010100001;
            14'h1f66: o_data_a = 16'b1110101010000111;
            14'h1f67: o_data_a = 16'b0000000000000001;
            14'h1f68: o_data_a = 16'b1111110111100000;
            14'h1f69: o_data_a = 16'b1110110111100000;
            14'h1f6a: o_data_a = 16'b1111110000010000;
            14'h1f6b: o_data_a = 16'b0000000000000000;
            14'h1f6c: o_data_a = 16'b1111110111101000;
            14'h1f6d: o_data_a = 16'b1110110010100000;
            14'h1f6e: o_data_a = 16'b1110001100001000;
            14'h1f6f: o_data_a = 16'b0000000000000000;
            14'h1f70: o_data_a = 16'b1111110010101000;
            14'h1f71: o_data_a = 16'b1111110000010000;
            14'h1f72: o_data_a = 16'b0001111101110110;
            14'h1f73: o_data_a = 16'b1110001100000101;
            14'h1f74: o_data_a = 16'b0001111110000111;
            14'h1f75: o_data_a = 16'b1110101010000111;
            14'h1f76: o_data_a = 16'b0000000000000001;
            14'h1f77: o_data_a = 16'b1111110111100000;
            14'h1f78: o_data_a = 16'b1111110000010000;
            14'h1f79: o_data_a = 16'b0000000000000000;
            14'h1f7a: o_data_a = 16'b1111110111101000;
            14'h1f7b: o_data_a = 16'b1110110010100000;
            14'h1f7c: o_data_a = 16'b1110001100001000;
            14'h1f7d: o_data_a = 16'b0000000000000000;
            14'h1f7e: o_data_a = 16'b1111110010100000;
            14'h1f7f: o_data_a = 16'b1111110001010000;
            14'h1f80: o_data_a = 16'b1110011111001000;
            14'h1f81: o_data_a = 16'b0000000000000000;
            14'h1f82: o_data_a = 16'b1111110010101000;
            14'h1f83: o_data_a = 16'b1111110000010000;
            14'h1f84: o_data_a = 16'b0000000000000001;
            14'h1f85: o_data_a = 16'b1111110111100000;
            14'h1f86: o_data_a = 16'b1110001100001000;
            14'h1f87: o_data_a = 16'b0000000000000001;
            14'h1f88: o_data_a = 16'b1111110111100000;
            14'h1f89: o_data_a = 16'b1111110000010000;
            14'h1f8a: o_data_a = 16'b0000000000000000;
            14'h1f8b: o_data_a = 16'b1111110111101000;
            14'h1f8c: o_data_a = 16'b1110110010100000;
            14'h1f8d: o_data_a = 16'b1110001100001000;
            14'h1f8e: o_data_a = 16'b0000000000110110;
            14'h1f8f: o_data_a = 16'b1110101010000111;
            14'h1f90: o_data_a = 16'b0000000000000100;
            14'h1f91: o_data_a = 16'b1110110000010000;
            14'h1f92: o_data_a = 16'b1110001110010000;
            14'h1f93: o_data_a = 16'b0000000000000000;
            14'h1f94: o_data_a = 16'b1111110111101000;
            14'h1f95: o_data_a = 16'b1110110010100000;
            14'h1f96: o_data_a = 16'b1110101010001000;
            14'h1f97: o_data_a = 16'b0001111110010010;
            14'h1f98: o_data_a = 16'b1110001100000001;
            14'h1f99: o_data_a = 16'b0000000000000010;
            14'h1f9a: o_data_a = 16'b1111110000100000;
            14'h1f9b: o_data_a = 16'b1111110000010000;
            14'h1f9c: o_data_a = 16'b0000000000000000;
            14'h1f9d: o_data_a = 16'b1111110111101000;
            14'h1f9e: o_data_a = 16'b1110110010100000;
            14'h1f9f: o_data_a = 16'b1110001100001000;
            14'h1fa0: o_data_a = 16'b0000000000000000;
            14'h1fa1: o_data_a = 16'b1111110111001000;
            14'h1fa2: o_data_a = 16'b1111110010100000;
            14'h1fa3: o_data_a = 16'b1110101010001000;
            14'h1fa4: o_data_a = 16'b0001111110101000;
            14'h1fa5: o_data_a = 16'b1110110000010000;
            14'h1fa6: o_data_a = 16'b0000000000100110;
            14'h1fa7: o_data_a = 16'b1110101010000111;
            14'h1fa8: o_data_a = 16'b0000000000000000;
            14'h1fa9: o_data_a = 16'b1111110010101000;
            14'h1faa: o_data_a = 16'b1111110000010000;
            14'h1fab: o_data_a = 16'b0001111110101111;
            14'h1fac: o_data_a = 16'b1110001100000101;
            14'h1fad: o_data_a = 16'b0001111111000110;
            14'h1fae: o_data_a = 16'b1110101010000111;
            14'h1faf: o_data_a = 16'b0000000000000100;
            14'h1fb0: o_data_a = 16'b1110110000010000;
            14'h1fb1: o_data_a = 16'b0000000000000000;
            14'h1fb2: o_data_a = 16'b1111110111101000;
            14'h1fb3: o_data_a = 16'b1110110010100000;
            14'h1fb4: o_data_a = 16'b1110001100001000;
            14'h1fb5: o_data_a = 16'b0000000000000001;
            14'h1fb6: o_data_a = 16'b1110110000010000;
            14'h1fb7: o_data_a = 16'b0000000000001101;
            14'h1fb8: o_data_a = 16'b1110001100001000;
            14'h1fb9: o_data_a = 16'b0110101011011001;
            14'h1fba: o_data_a = 16'b1110110000010000;
            14'h1fbb: o_data_a = 16'b0000000000001110;
            14'h1fbc: o_data_a = 16'b1110001100001000;
            14'h1fbd: o_data_a = 16'b0001111111000001;
            14'h1fbe: o_data_a = 16'b1110110000010000;
            14'h1fbf: o_data_a = 16'b0000000001011111;
            14'h1fc0: o_data_a = 16'b1110101010000111;
            14'h1fc1: o_data_a = 16'b0000000000000000;
            14'h1fc2: o_data_a = 16'b1111110010101000;
            14'h1fc3: o_data_a = 16'b1111110000010000;
            14'h1fc4: o_data_a = 16'b0000000000000101;
            14'h1fc5: o_data_a = 16'b1110001100001000;
            14'h1fc6: o_data_a = 16'b0000000000000111;
            14'h1fc7: o_data_a = 16'b1110110000010000;
            14'h1fc8: o_data_a = 16'b0000000000000000;
            14'h1fc9: o_data_a = 16'b1111110111101000;
            14'h1fca: o_data_a = 16'b1110110010100000;
            14'h1fcb: o_data_a = 16'b1110001100001000;
            14'h1fcc: o_data_a = 16'b0000000000000000;
            14'h1fcd: o_data_a = 16'b1111110010101000;
            14'h1fce: o_data_a = 16'b1111110000010000;
            14'h1fcf: o_data_a = 16'b0000000000000001;
            14'h1fd0: o_data_a = 16'b1111110000100000;
            14'h1fd1: o_data_a = 16'b1110001100001000;
            14'h1fd2: o_data_a = 16'b0000000000000001;
            14'h1fd3: o_data_a = 16'b1111110000100000;
            14'h1fd4: o_data_a = 16'b1111110000010000;
            14'h1fd5: o_data_a = 16'b0000000000000000;
            14'h1fd6: o_data_a = 16'b1111110111101000;
            14'h1fd7: o_data_a = 16'b1110110010100000;
            14'h1fd8: o_data_a = 16'b1110001100001000;
            14'h1fd9: o_data_a = 16'b0000000000000000;
            14'h1fda: o_data_a = 16'b1111110111001000;
            14'h1fdb: o_data_a = 16'b1111110010100000;
            14'h1fdc: o_data_a = 16'b1110111111001000;
            14'h1fdd: o_data_a = 16'b0000000000000000;
            14'h1fde: o_data_a = 16'b1111110010100000;
            14'h1fdf: o_data_a = 16'b1111110001010000;
            14'h1fe0: o_data_a = 16'b1110011111001000;
            14'h1fe1: o_data_a = 16'b0001111111100101;
            14'h1fe2: o_data_a = 16'b1110110000010000;
            14'h1fe3: o_data_a = 16'b0000000000010110;
            14'h1fe4: o_data_a = 16'b1110101010000111;
            14'h1fe5: o_data_a = 16'b0000000000000000;
            14'h1fe6: o_data_a = 16'b1111110010100000;
            14'h1fe7: o_data_a = 16'b1111110001001000;
            14'h1fe8: o_data_a = 16'b0000000000000000;
            14'h1fe9: o_data_a = 16'b1111110010101000;
            14'h1fea: o_data_a = 16'b1111110000010000;
            14'h1feb: o_data_a = 16'b0010000010011100;
            14'h1fec: o_data_a = 16'b1110001100000101;
            14'h1fed: o_data_a = 16'b0000000000000001;
            14'h1fee: o_data_a = 16'b1111110000010000;
            14'h1fef: o_data_a = 16'b0000000000000011;
            14'h1ff0: o_data_a = 16'b1110000010100000;
            14'h1ff1: o_data_a = 16'b1111110000010000;
            14'h1ff2: o_data_a = 16'b0000000000000000;
            14'h1ff3: o_data_a = 16'b1111110111101000;
            14'h1ff4: o_data_a = 16'b1110110010100000;
            14'h1ff5: o_data_a = 16'b1110001100001000;
            14'h1ff6: o_data_a = 16'b0000000000000001;
            14'h1ff7: o_data_a = 16'b1111110000100000;
            14'h1ff8: o_data_a = 16'b1111110000010000;
            14'h1ff9: o_data_a = 16'b0000000000000000;
            14'h1ffa: o_data_a = 16'b1111110111101000;
            14'h1ffb: o_data_a = 16'b1110110010100000;
            14'h1ffc: o_data_a = 16'b1110001100001000;
            14'h1ffd: o_data_a = 16'b0000000000010010;
            14'h1ffe: o_data_a = 16'b1111110000010000;
            14'h1fff: o_data_a = 16'b0000000000000000;
            14'h2000: o_data_a = 16'b1111110111101000;
            14'h2001: o_data_a = 16'b1110110010100000;
            14'h2002: o_data_a = 16'b1110001100001000;
            14'h2003: o_data_a = 16'b0000000000000000;
            14'h2004: o_data_a = 16'b1111110010101000;
            14'h2005: o_data_a = 16'b1111110000010000;
            14'h2006: o_data_a = 16'b1110110010100000;
            14'h2007: o_data_a = 16'b1111000010001000;
            14'h2008: o_data_a = 16'b0000000000000000;
            14'h2009: o_data_a = 16'b1111110010101000;
            14'h200a: o_data_a = 16'b1111110000010000;
            14'h200b: o_data_a = 16'b0000000000000100;
            14'h200c: o_data_a = 16'b1110001100001000;
            14'h200d: o_data_a = 16'b0000000000000100;
            14'h200e: o_data_a = 16'b1111110000100000;
            14'h200f: o_data_a = 16'b1111110000010000;
            14'h2010: o_data_a = 16'b0000000000000000;
            14'h2011: o_data_a = 16'b1111110111101000;
            14'h2012: o_data_a = 16'b1110110010100000;
            14'h2013: o_data_a = 16'b1110001100001000;
            14'h2014: o_data_a = 16'b0000000000000000;
            14'h2015: o_data_a = 16'b1111110010101000;
            14'h2016: o_data_a = 16'b1111110000010000;
            14'h2017: o_data_a = 16'b1110110010100000;
            14'h2018: o_data_a = 16'b1111000010001000;
            14'h2019: o_data_a = 16'b0000000000000000;
            14'h201a: o_data_a = 16'b1111110010101000;
            14'h201b: o_data_a = 16'b1111110000010000;
            14'h201c: o_data_a = 16'b0000000000000001;
            14'h201d: o_data_a = 16'b1111110111100000;
            14'h201e: o_data_a = 16'b1110001100001000;
            14'h201f: o_data_a = 16'b0000000000000001;
            14'h2020: o_data_a = 16'b1111110111100000;
            14'h2021: o_data_a = 16'b1111110000010000;
            14'h2022: o_data_a = 16'b0000000000000000;
            14'h2023: o_data_a = 16'b1111110111101000;
            14'h2024: o_data_a = 16'b1110110010100000;
            14'h2025: o_data_a = 16'b1110001100001000;
            14'h2026: o_data_a = 16'b0000000000000001;
            14'h2027: o_data_a = 16'b1111110111100000;
            14'h2028: o_data_a = 16'b1111110000010000;
            14'h2029: o_data_a = 16'b0000000000000000;
            14'h202a: o_data_a = 16'b1111110111101000;
            14'h202b: o_data_a = 16'b1110110010100000;
            14'h202c: o_data_a = 16'b1110001100001000;
            14'h202d: o_data_a = 16'b0000000000000010;
            14'h202e: o_data_a = 16'b1110110000010000;
            14'h202f: o_data_a = 16'b0000000000001101;
            14'h2030: o_data_a = 16'b1110001100001000;
            14'h2031: o_data_a = 16'b0001101010100110;
            14'h2032: o_data_a = 16'b1110110000010000;
            14'h2033: o_data_a = 16'b0000000000001110;
            14'h2034: o_data_a = 16'b1110001100001000;
            14'h2035: o_data_a = 16'b0010000000111001;
            14'h2036: o_data_a = 16'b1110110000010000;
            14'h2037: o_data_a = 16'b0000000001011111;
            14'h2038: o_data_a = 16'b1110101010000111;
            14'h2039: o_data_a = 16'b0000000000000000;
            14'h203a: o_data_a = 16'b1111110010101000;
            14'h203b: o_data_a = 16'b1111110000010000;
            14'h203c: o_data_a = 16'b0000000000000001;
            14'h203d: o_data_a = 16'b1111110111100000;
            14'h203e: o_data_a = 16'b1110110111100000;
            14'h203f: o_data_a = 16'b1110001100001000;
            14'h2040: o_data_a = 16'b0000000000000001;
            14'h2041: o_data_a = 16'b1111110111100000;
            14'h2042: o_data_a = 16'b1110110111100000;
            14'h2043: o_data_a = 16'b1111110000010000;
            14'h2044: o_data_a = 16'b0000000000000000;
            14'h2045: o_data_a = 16'b1111110111101000;
            14'h2046: o_data_a = 16'b1110110010100000;
            14'h2047: o_data_a = 16'b1110001100001000;
            14'h2048: o_data_a = 16'b0000000000000010;
            14'h2049: o_data_a = 16'b1111110000100000;
            14'h204a: o_data_a = 16'b1111110000010000;
            14'h204b: o_data_a = 16'b0000000000000000;
            14'h204c: o_data_a = 16'b1111110111101000;
            14'h204d: o_data_a = 16'b1110110010100000;
            14'h204e: o_data_a = 16'b1110001100001000;
            14'h204f: o_data_a = 16'b0010000001010011;
            14'h2050: o_data_a = 16'b1110110000010000;
            14'h2051: o_data_a = 16'b0000000000010110;
            14'h2052: o_data_a = 16'b1110101010000111;
            14'h2053: o_data_a = 16'b0000000000000000;
            14'h2054: o_data_a = 16'b1111110010100000;
            14'h2055: o_data_a = 16'b1111110001001000;
            14'h2056: o_data_a = 16'b0000000000000001;
            14'h2057: o_data_a = 16'b1111110111100000;
            14'h2058: o_data_a = 16'b1110110111100000;
            14'h2059: o_data_a = 16'b1111110000010000;
            14'h205a: o_data_a = 16'b0000000000000000;
            14'h205b: o_data_a = 16'b1111110111101000;
            14'h205c: o_data_a = 16'b1110110010100000;
            14'h205d: o_data_a = 16'b1110001100001000;
            14'h205e: o_data_a = 16'b0000000000000000;
            14'h205f: o_data_a = 16'b1111110111001000;
            14'h2060: o_data_a = 16'b1111110010100000;
            14'h2061: o_data_a = 16'b1110101010001000;
            14'h2062: o_data_a = 16'b0010000001100110;
            14'h2063: o_data_a = 16'b1110110000010000;
            14'h2064: o_data_a = 16'b0000000000100110;
            14'h2065: o_data_a = 16'b1110101010000111;
            14'h2066: o_data_a = 16'b0000000000000000;
            14'h2067: o_data_a = 16'b1111110010100000;
            14'h2068: o_data_a = 16'b1111110001001000;
            14'h2069: o_data_a = 16'b0000000000000000;
            14'h206a: o_data_a = 16'b1111110010101000;
            14'h206b: o_data_a = 16'b1111110000010000;
            14'h206c: o_data_a = 16'b1110110010100000;
            14'h206d: o_data_a = 16'b1111000000001000;
            14'h206e: o_data_a = 16'b0000000000000000;
            14'h206f: o_data_a = 16'b1111110010101000;
            14'h2070: o_data_a = 16'b1111110000010000;
            14'h2071: o_data_a = 16'b0010000001110101;
            14'h2072: o_data_a = 16'b1110001100000101;
            14'h2073: o_data_a = 16'b0010000010000100;
            14'h2074: o_data_a = 16'b1110101010000111;
            14'h2075: o_data_a = 16'b0000000000000001;
            14'h2076: o_data_a = 16'b1111110111100000;
            14'h2077: o_data_a = 16'b1111110000010000;
            14'h2078: o_data_a = 16'b0000000000000000;
            14'h2079: o_data_a = 16'b1111110111101000;
            14'h207a: o_data_a = 16'b1110110010100000;
            14'h207b: o_data_a = 16'b1110001100001000;
            14'h207c: o_data_a = 16'b0000000000000000;
            14'h207d: o_data_a = 16'b1111110010101000;
            14'h207e: o_data_a = 16'b1111110000010000;
            14'h207f: o_data_a = 16'b0000000000000001;
            14'h2080: o_data_a = 16'b1111110111100000;
            14'h2081: o_data_a = 16'b1110110111100000;
            14'h2082: o_data_a = 16'b1110110111100000;
            14'h2083: o_data_a = 16'b1110001100001000;
            14'h2084: o_data_a = 16'b0000000000000001;
            14'h2085: o_data_a = 16'b1111110000100000;
            14'h2086: o_data_a = 16'b1111110000010000;
            14'h2087: o_data_a = 16'b0000000000000000;
            14'h2088: o_data_a = 16'b1111110111101000;
            14'h2089: o_data_a = 16'b1110110010100000;
            14'h208a: o_data_a = 16'b1110001100001000;
            14'h208b: o_data_a = 16'b0000000000000000;
            14'h208c: o_data_a = 16'b1111110111001000;
            14'h208d: o_data_a = 16'b1111110010100000;
            14'h208e: o_data_a = 16'b1110111111001000;
            14'h208f: o_data_a = 16'b0000000000000000;
            14'h2090: o_data_a = 16'b1111110010101000;
            14'h2091: o_data_a = 16'b1111110000010000;
            14'h2092: o_data_a = 16'b1110110010100000;
            14'h2093: o_data_a = 16'b1111000111001000;
            14'h2094: o_data_a = 16'b0000000000000000;
            14'h2095: o_data_a = 16'b1111110010101000;
            14'h2096: o_data_a = 16'b1111110000010000;
            14'h2097: o_data_a = 16'b0000000000000001;
            14'h2098: o_data_a = 16'b1111110000100000;
            14'h2099: o_data_a = 16'b1110001100001000;
            14'h209a: o_data_a = 16'b0001111111010010;
            14'h209b: o_data_a = 16'b1110101010000111;
            14'h209c: o_data_a = 16'b0000000000000001;
            14'h209d: o_data_a = 16'b1111110000010000;
            14'h209e: o_data_a = 16'b0000000000000011;
            14'h209f: o_data_a = 16'b1110000010100000;
            14'h20a0: o_data_a = 16'b1111110000010000;
            14'h20a1: o_data_a = 16'b0000000000000000;
            14'h20a2: o_data_a = 16'b1111110111101000;
            14'h20a3: o_data_a = 16'b1110110010100000;
            14'h20a4: o_data_a = 16'b1110001100001000;
            14'h20a5: o_data_a = 16'b0000000000110110;
            14'h20a6: o_data_a = 16'b1110101010000111;
            14'h20a7: o_data_a = 16'b0000000000000010;
            14'h20a8: o_data_a = 16'b1111110000100000;
            14'h20a9: o_data_a = 16'b1111110000010000;
            14'h20aa: o_data_a = 16'b0000000000000000;
            14'h20ab: o_data_a = 16'b1111110111101000;
            14'h20ac: o_data_a = 16'b1110110010100000;
            14'h20ad: o_data_a = 16'b1110001100001000;
            14'h20ae: o_data_a = 16'b0000000000000010;
            14'h20af: o_data_a = 16'b1111110111100000;
            14'h20b0: o_data_a = 16'b1111110000010000;
            14'h20b1: o_data_a = 16'b0000000000000000;
            14'h20b2: o_data_a = 16'b1111110111101000;
            14'h20b3: o_data_a = 16'b1110110010100000;
            14'h20b4: o_data_a = 16'b1110001100001000;
            14'h20b5: o_data_a = 16'b0010000010111001;
            14'h20b6: o_data_a = 16'b1110110000010000;
            14'h20b7: o_data_a = 16'b0000000000010110;
            14'h20b8: o_data_a = 16'b1110101010000111;
            14'h20b9: o_data_a = 16'b0000000000000000;
            14'h20ba: o_data_a = 16'b1111110010101000;
            14'h20bb: o_data_a = 16'b1111110000010000;
            14'h20bc: o_data_a = 16'b0010000011000000;
            14'h20bd: o_data_a = 16'b1110001100000101;
            14'h20be: o_data_a = 16'b0010000011001101;
            14'h20bf: o_data_a = 16'b1110101010000111;
            14'h20c0: o_data_a = 16'b0000000000000010;
            14'h20c1: o_data_a = 16'b1111110000100000;
            14'h20c2: o_data_a = 16'b1111110000010000;
            14'h20c3: o_data_a = 16'b0000000000000000;
            14'h20c4: o_data_a = 16'b1111110111101000;
            14'h20c5: o_data_a = 16'b1110110010100000;
            14'h20c6: o_data_a = 16'b1110001100001000;
            14'h20c7: o_data_a = 16'b0000000000000000;
            14'h20c8: o_data_a = 16'b1111110010101000;
            14'h20c9: o_data_a = 16'b1111110000010000;
            14'h20ca: o_data_a = 16'b0000000000000010;
            14'h20cb: o_data_a = 16'b1111110111100000;
            14'h20cc: o_data_a = 16'b1110001100001000;
            14'h20cd: o_data_a = 16'b0000000000000010;
            14'h20ce: o_data_a = 16'b1111110111100000;
            14'h20cf: o_data_a = 16'b1111110000010000;
            14'h20d0: o_data_a = 16'b0000000000000000;
            14'h20d1: o_data_a = 16'b1111110111101000;
            14'h20d2: o_data_a = 16'b1110110010100000;
            14'h20d3: o_data_a = 16'b1110001100001000;
            14'h20d4: o_data_a = 16'b0000000000110110;
            14'h20d5: o_data_a = 16'b1110101010000111;
            14'h20d6: o_data_a = 16'b0000000000000010;
            14'h20d7: o_data_a = 16'b1111110000100000;
            14'h20d8: o_data_a = 16'b1111110000010000;
            14'h20d9: o_data_a = 16'b0000000000000000;
            14'h20da: o_data_a = 16'b1111110111101000;
            14'h20db: o_data_a = 16'b1110110010100000;
            14'h20dc: o_data_a = 16'b1110001100001000;
            14'h20dd: o_data_a = 16'b0000000000000010;
            14'h20de: o_data_a = 16'b1111110111100000;
            14'h20df: o_data_a = 16'b1111110000010000;
            14'h20e0: o_data_a = 16'b0000000000000000;
            14'h20e1: o_data_a = 16'b1111110111101000;
            14'h20e2: o_data_a = 16'b1110110010100000;
            14'h20e3: o_data_a = 16'b1110001100001000;
            14'h20e4: o_data_a = 16'b0010000011101000;
            14'h20e5: o_data_a = 16'b1110110000010000;
            14'h20e6: o_data_a = 16'b0000000000100110;
            14'h20e7: o_data_a = 16'b1110101010000111;
            14'h20e8: o_data_a = 16'b0000000000000000;
            14'h20e9: o_data_a = 16'b1111110010101000;
            14'h20ea: o_data_a = 16'b1111110000010000;
            14'h20eb: o_data_a = 16'b0010000011101111;
            14'h20ec: o_data_a = 16'b1110001100000101;
            14'h20ed: o_data_a = 16'b0010000011111100;
            14'h20ee: o_data_a = 16'b1110101010000111;
            14'h20ef: o_data_a = 16'b0000000000000010;
            14'h20f0: o_data_a = 16'b1111110000100000;
            14'h20f1: o_data_a = 16'b1111110000010000;
            14'h20f2: o_data_a = 16'b0000000000000000;
            14'h20f3: o_data_a = 16'b1111110111101000;
            14'h20f4: o_data_a = 16'b1110110010100000;
            14'h20f5: o_data_a = 16'b1110001100001000;
            14'h20f6: o_data_a = 16'b0000000000000000;
            14'h20f7: o_data_a = 16'b1111110010101000;
            14'h20f8: o_data_a = 16'b1111110000010000;
            14'h20f9: o_data_a = 16'b0000000000000010;
            14'h20fa: o_data_a = 16'b1111110111100000;
            14'h20fb: o_data_a = 16'b1110001100001000;
            14'h20fc: o_data_a = 16'b0000000000000010;
            14'h20fd: o_data_a = 16'b1111110111100000;
            14'h20fe: o_data_a = 16'b1111110000010000;
            14'h20ff: o_data_a = 16'b0000000000000000;
            14'h2100: o_data_a = 16'b1111110111101000;
            14'h2101: o_data_a = 16'b1110110010100000;
            14'h2102: o_data_a = 16'b1110001100001000;
            14'h2103: o_data_a = 16'b0000000000110110;
            14'h2104: o_data_a = 16'b1110101010000111;
            14'h2105: o_data_a = 16'b0000000000000000;
            14'h2106: o_data_a = 16'b1111110111001000;
            14'h2107: o_data_a = 16'b1111110010100000;
            14'h2108: o_data_a = 16'b1110101010001000;
            14'h2109: o_data_a = 16'b0000000000000000;
            14'h210a: o_data_a = 16'b1111110010101000;
            14'h210b: o_data_a = 16'b1111110000010000;
            14'h210c: o_data_a = 16'b0000000000010011;
            14'h210d: o_data_a = 16'b1110001100001000;
            14'h210e: o_data_a = 16'b0000100000000000;
            14'h210f: o_data_a = 16'b1110110000010000;
            14'h2110: o_data_a = 16'b0000000000000000;
            14'h2111: o_data_a = 16'b1111110111101000;
            14'h2112: o_data_a = 16'b1110110010100000;
            14'h2113: o_data_a = 16'b1110001100001000;
            14'h2114: o_data_a = 16'b0000000000010011;
            14'h2115: o_data_a = 16'b1111110000010000;
            14'h2116: o_data_a = 16'b0000000000000000;
            14'h2117: o_data_a = 16'b1111110111101000;
            14'h2118: o_data_a = 16'b1110110010100000;
            14'h2119: o_data_a = 16'b1110001100001000;
            14'h211a: o_data_a = 16'b0000000000000000;
            14'h211b: o_data_a = 16'b1111110010101000;
            14'h211c: o_data_a = 16'b1111110000010000;
            14'h211d: o_data_a = 16'b1110110010100000;
            14'h211e: o_data_a = 16'b1111000010001000;
            14'h211f: o_data_a = 16'b0011011111111110;
            14'h2120: o_data_a = 16'b1110110000010000;
            14'h2121: o_data_a = 16'b0000000000000000;
            14'h2122: o_data_a = 16'b1111110111101000;
            14'h2123: o_data_a = 16'b1110110010100000;
            14'h2124: o_data_a = 16'b1110001100001000;
            14'h2125: o_data_a = 16'b0000000000000000;
            14'h2126: o_data_a = 16'b1111110010101000;
            14'h2127: o_data_a = 16'b1111110000010000;
            14'h2128: o_data_a = 16'b0000000000000101;
            14'h2129: o_data_a = 16'b1110001100001000;
            14'h212a: o_data_a = 16'b0000000000000000;
            14'h212b: o_data_a = 16'b1111110010101000;
            14'h212c: o_data_a = 16'b1111110000010000;
            14'h212d: o_data_a = 16'b0000000000000100;
            14'h212e: o_data_a = 16'b1110001100001000;
            14'h212f: o_data_a = 16'b0000000000000101;
            14'h2130: o_data_a = 16'b1111110000010000;
            14'h2131: o_data_a = 16'b0000000000000000;
            14'h2132: o_data_a = 16'b1111110111101000;
            14'h2133: o_data_a = 16'b1110110010100000;
            14'h2134: o_data_a = 16'b1110001100001000;
            14'h2135: o_data_a = 16'b0000000000000000;
            14'h2136: o_data_a = 16'b1111110010101000;
            14'h2137: o_data_a = 16'b1111110000010000;
            14'h2138: o_data_a = 16'b0000000000000100;
            14'h2139: o_data_a = 16'b1111110000100000;
            14'h213a: o_data_a = 16'b1110001100001000;
            14'h213b: o_data_a = 16'b0000100000000001;
            14'h213c: o_data_a = 16'b1110110000010000;
            14'h213d: o_data_a = 16'b0000000000000000;
            14'h213e: o_data_a = 16'b1111110111101000;
            14'h213f: o_data_a = 16'b1110110010100000;
            14'h2140: o_data_a = 16'b1110001100001000;
            14'h2141: o_data_a = 16'b0000000000010011;
            14'h2142: o_data_a = 16'b1111110000010000;
            14'h2143: o_data_a = 16'b0000000000000000;
            14'h2144: o_data_a = 16'b1111110111101000;
            14'h2145: o_data_a = 16'b1110110010100000;
            14'h2146: o_data_a = 16'b1110001100001000;
            14'h2147: o_data_a = 16'b0000000000000000;
            14'h2148: o_data_a = 16'b1111110010101000;
            14'h2149: o_data_a = 16'b1111110000010000;
            14'h214a: o_data_a = 16'b1110110010100000;
            14'h214b: o_data_a = 16'b1111000010001000;
            14'h214c: o_data_a = 16'b0000100000000010;
            14'h214d: o_data_a = 16'b1110110000010000;
            14'h214e: o_data_a = 16'b0000000000000000;
            14'h214f: o_data_a = 16'b1111110111101000;
            14'h2150: o_data_a = 16'b1110110010100000;
            14'h2151: o_data_a = 16'b1110001100001000;
            14'h2152: o_data_a = 16'b0000000000000000;
            14'h2153: o_data_a = 16'b1111110010101000;
            14'h2154: o_data_a = 16'b1111110000010000;
            14'h2155: o_data_a = 16'b0000000000000101;
            14'h2156: o_data_a = 16'b1110001100001000;
            14'h2157: o_data_a = 16'b0000000000000000;
            14'h2158: o_data_a = 16'b1111110010101000;
            14'h2159: o_data_a = 16'b1111110000010000;
            14'h215a: o_data_a = 16'b0000000000000100;
            14'h215b: o_data_a = 16'b1110001100001000;
            14'h215c: o_data_a = 16'b0000000000000101;
            14'h215d: o_data_a = 16'b1111110000010000;
            14'h215e: o_data_a = 16'b0000000000000000;
            14'h215f: o_data_a = 16'b1111110111101000;
            14'h2160: o_data_a = 16'b1110110010100000;
            14'h2161: o_data_a = 16'b1110001100001000;
            14'h2162: o_data_a = 16'b0000000000000000;
            14'h2163: o_data_a = 16'b1111110010101000;
            14'h2164: o_data_a = 16'b1111110000010000;
            14'h2165: o_data_a = 16'b0000000000000100;
            14'h2166: o_data_a = 16'b1111110000100000;
            14'h2167: o_data_a = 16'b1110001100001000;
            14'h2168: o_data_a = 16'b0000000000000000;
            14'h2169: o_data_a = 16'b1111110111001000;
            14'h216a: o_data_a = 16'b1111110010100000;
            14'h216b: o_data_a = 16'b1110101010001000;
            14'h216c: o_data_a = 16'b0000000000110110;
            14'h216d: o_data_a = 16'b1110101010000111;
            14'h216e: o_data_a = 16'b0000000000000010;
            14'h216f: o_data_a = 16'b1111110000100000;
            14'h2170: o_data_a = 16'b1111110000010000;
            14'h2171: o_data_a = 16'b0000000000000000;
            14'h2172: o_data_a = 16'b1111110111101000;
            14'h2173: o_data_a = 16'b1110110010100000;
            14'h2174: o_data_a = 16'b1110001100001000;
            14'h2175: o_data_a = 16'b0000000000010011;
            14'h2176: o_data_a = 16'b1111110000010000;
            14'h2177: o_data_a = 16'b0000000000000000;
            14'h2178: o_data_a = 16'b1111110111101000;
            14'h2179: o_data_a = 16'b1110110010100000;
            14'h217a: o_data_a = 16'b1110001100001000;
            14'h217b: o_data_a = 16'b0000000000000000;
            14'h217c: o_data_a = 16'b1111110010101000;
            14'h217d: o_data_a = 16'b1111110000010000;
            14'h217e: o_data_a = 16'b1110110010100000;
            14'h217f: o_data_a = 16'b1111000010001000;
            14'h2180: o_data_a = 16'b0000000000000000;
            14'h2181: o_data_a = 16'b1111110010101000;
            14'h2182: o_data_a = 16'b1111110000010000;
            14'h2183: o_data_a = 16'b0000000000000100;
            14'h2184: o_data_a = 16'b1110001100001000;
            14'h2185: o_data_a = 16'b0000000000000100;
            14'h2186: o_data_a = 16'b1111110000100000;
            14'h2187: o_data_a = 16'b1111110000010000;
            14'h2188: o_data_a = 16'b0000000000000000;
            14'h2189: o_data_a = 16'b1111110111101000;
            14'h218a: o_data_a = 16'b1110110010100000;
            14'h218b: o_data_a = 16'b1110001100001000;
            14'h218c: o_data_a = 16'b0000000000110110;
            14'h218d: o_data_a = 16'b1110101010000111;
            14'h218e: o_data_a = 16'b0000000000000010;
            14'h218f: o_data_a = 16'b1111110000100000;
            14'h2190: o_data_a = 16'b1111110000010000;
            14'h2191: o_data_a = 16'b0000000000000000;
            14'h2192: o_data_a = 16'b1111110111101000;
            14'h2193: o_data_a = 16'b1110110010100000;
            14'h2194: o_data_a = 16'b1110001100001000;
            14'h2195: o_data_a = 16'b0000000000010011;
            14'h2196: o_data_a = 16'b1111110000010000;
            14'h2197: o_data_a = 16'b0000000000000000;
            14'h2198: o_data_a = 16'b1111110111101000;
            14'h2199: o_data_a = 16'b1110110010100000;
            14'h219a: o_data_a = 16'b1110001100001000;
            14'h219b: o_data_a = 16'b0000000000000000;
            14'h219c: o_data_a = 16'b1111110010101000;
            14'h219d: o_data_a = 16'b1111110000010000;
            14'h219e: o_data_a = 16'b1110110010100000;
            14'h219f: o_data_a = 16'b1111000010001000;
            14'h21a0: o_data_a = 16'b0000000000000010;
            14'h21a1: o_data_a = 16'b1111110111100000;
            14'h21a2: o_data_a = 16'b1111110000010000;
            14'h21a3: o_data_a = 16'b0000000000000000;
            14'h21a4: o_data_a = 16'b1111110111101000;
            14'h21a5: o_data_a = 16'b1110110010100000;
            14'h21a6: o_data_a = 16'b1110001100001000;
            14'h21a7: o_data_a = 16'b0000000000000000;
            14'h21a8: o_data_a = 16'b1111110010101000;
            14'h21a9: o_data_a = 16'b1111110000010000;
            14'h21aa: o_data_a = 16'b0000000000000101;
            14'h21ab: o_data_a = 16'b1110001100001000;
            14'h21ac: o_data_a = 16'b0000000000000000;
            14'h21ad: o_data_a = 16'b1111110010101000;
            14'h21ae: o_data_a = 16'b1111110000010000;
            14'h21af: o_data_a = 16'b0000000000000100;
            14'h21b0: o_data_a = 16'b1110001100001000;
            14'h21b1: o_data_a = 16'b0000000000000101;
            14'h21b2: o_data_a = 16'b1111110000010000;
            14'h21b3: o_data_a = 16'b0000000000000000;
            14'h21b4: o_data_a = 16'b1111110111101000;
            14'h21b5: o_data_a = 16'b1110110010100000;
            14'h21b6: o_data_a = 16'b1110001100001000;
            14'h21b7: o_data_a = 16'b0000000000000000;
            14'h21b8: o_data_a = 16'b1111110010101000;
            14'h21b9: o_data_a = 16'b1111110000010000;
            14'h21ba: o_data_a = 16'b0000000000000100;
            14'h21bb: o_data_a = 16'b1111110000100000;
            14'h21bc: o_data_a = 16'b1110001100001000;
            14'h21bd: o_data_a = 16'b0000000000000000;
            14'h21be: o_data_a = 16'b1111110111001000;
            14'h21bf: o_data_a = 16'b1111110010100000;
            14'h21c0: o_data_a = 16'b1110101010001000;
            14'h21c1: o_data_a = 16'b0000000000110110;
            14'h21c2: o_data_a = 16'b1110101010000111;
            14'h21c3: o_data_a = 16'b0000000000000000;
            14'h21c4: o_data_a = 16'b1111110111101000;
            14'h21c5: o_data_a = 16'b1110110010100000;
            14'h21c6: o_data_a = 16'b1110101010001000;
            14'h21c7: o_data_a = 16'b0000000000000010;
            14'h21c8: o_data_a = 16'b1111110000100000;
            14'h21c9: o_data_a = 16'b1111110000010000;
            14'h21ca: o_data_a = 16'b0000000000000000;
            14'h21cb: o_data_a = 16'b1111110111101000;
            14'h21cc: o_data_a = 16'b1110110010100000;
            14'h21cd: o_data_a = 16'b1110001100001000;
            14'h21ce: o_data_a = 16'b0000000000000000;
            14'h21cf: o_data_a = 16'b1111110111001000;
            14'h21d0: o_data_a = 16'b1111110010100000;
            14'h21d1: o_data_a = 16'b1110111111001000;
            14'h21d2: o_data_a = 16'b0010000111010110;
            14'h21d3: o_data_a = 16'b1110110000010000;
            14'h21d4: o_data_a = 16'b0000000000100110;
            14'h21d5: o_data_a = 16'b1110101010000111;
            14'h21d6: o_data_a = 16'b0000000000000000;
            14'h21d7: o_data_a = 16'b1111110010101000;
            14'h21d8: o_data_a = 16'b1111110000010000;
            14'h21d9: o_data_a = 16'b0010000111011101;
            14'h21da: o_data_a = 16'b1110001100000101;
            14'h21db: o_data_a = 16'b0010000111110100;
            14'h21dc: o_data_a = 16'b1110101010000111;
            14'h21dd: o_data_a = 16'b0000000000000101;
            14'h21de: o_data_a = 16'b1110110000010000;
            14'h21df: o_data_a = 16'b0000000000000000;
            14'h21e0: o_data_a = 16'b1111110111101000;
            14'h21e1: o_data_a = 16'b1110110010100000;
            14'h21e2: o_data_a = 16'b1110001100001000;
            14'h21e3: o_data_a = 16'b0000000000000001;
            14'h21e4: o_data_a = 16'b1110110000010000;
            14'h21e5: o_data_a = 16'b0000000000001101;
            14'h21e6: o_data_a = 16'b1110001100001000;
            14'h21e7: o_data_a = 16'b0110101011011001;
            14'h21e8: o_data_a = 16'b1110110000010000;
            14'h21e9: o_data_a = 16'b0000000000001110;
            14'h21ea: o_data_a = 16'b1110001100001000;
            14'h21eb: o_data_a = 16'b0010000111101111;
            14'h21ec: o_data_a = 16'b1110110000010000;
            14'h21ed: o_data_a = 16'b0000000001011111;
            14'h21ee: o_data_a = 16'b1110101010000111;
            14'h21ef: o_data_a = 16'b0000000000000000;
            14'h21f0: o_data_a = 16'b1111110010101000;
            14'h21f1: o_data_a = 16'b1111110000010000;
            14'h21f2: o_data_a = 16'b0000000000000101;
            14'h21f3: o_data_a = 16'b1110001100001000;
            14'h21f4: o_data_a = 16'b0000100000000000;
            14'h21f5: o_data_a = 16'b1110110000010000;
            14'h21f6: o_data_a = 16'b0000000000000000;
            14'h21f7: o_data_a = 16'b1111110111101000;
            14'h21f8: o_data_a = 16'b1110110010100000;
            14'h21f9: o_data_a = 16'b1110001100001000;
            14'h21fa: o_data_a = 16'b0000000000000000;
            14'h21fb: o_data_a = 16'b1111110010101000;
            14'h21fc: o_data_a = 16'b1111110000010000;
            14'h21fd: o_data_a = 16'b0000000000000001;
            14'h21fe: o_data_a = 16'b1111110000100000;
            14'h21ff: o_data_a = 16'b1110001100001000;
            14'h2200: o_data_a = 16'b0000000000000000;
            14'h2201: o_data_a = 16'b1111110111001000;
            14'h2202: o_data_a = 16'b1111110010100000;
            14'h2203: o_data_a = 16'b1110101010001000;
            14'h2204: o_data_a = 16'b0000000000000001;
            14'h2205: o_data_a = 16'b1111110000100000;
            14'h2206: o_data_a = 16'b1111110000010000;
            14'h2207: o_data_a = 16'b0000000000000000;
            14'h2208: o_data_a = 16'b1111110111101000;
            14'h2209: o_data_a = 16'b1110110010100000;
            14'h220a: o_data_a = 16'b1110001100001000;
            14'h220b: o_data_a = 16'b0000000000000000;
            14'h220c: o_data_a = 16'b1111110010101000;
            14'h220d: o_data_a = 16'b1111110000010000;
            14'h220e: o_data_a = 16'b1110110010100000;
            14'h220f: o_data_a = 16'b1111000010001000;
            14'h2210: o_data_a = 16'b0000000000000000;
            14'h2211: o_data_a = 16'b1111110010101000;
            14'h2212: o_data_a = 16'b1111110000010000;
            14'h2213: o_data_a = 16'b0000000000000100;
            14'h2214: o_data_a = 16'b1110001100001000;
            14'h2215: o_data_a = 16'b0000000000000100;
            14'h2216: o_data_a = 16'b1111110000100000;
            14'h2217: o_data_a = 16'b1111110000010000;
            14'h2218: o_data_a = 16'b0000000000000000;
            14'h2219: o_data_a = 16'b1111110111101000;
            14'h221a: o_data_a = 16'b1110110010100000;
            14'h221b: o_data_a = 16'b1110001100001000;
            14'h221c: o_data_a = 16'b0000000000000010;
            14'h221d: o_data_a = 16'b1111110000100000;
            14'h221e: o_data_a = 16'b1111110000010000;
            14'h221f: o_data_a = 16'b0000000000000000;
            14'h2220: o_data_a = 16'b1111110111101000;
            14'h2221: o_data_a = 16'b1110110010100000;
            14'h2222: o_data_a = 16'b1110001100001000;
            14'h2223: o_data_a = 16'b0010001000100111;
            14'h2224: o_data_a = 16'b1110110000010000;
            14'h2225: o_data_a = 16'b0000000000100110;
            14'h2226: o_data_a = 16'b1110101010000111;
            14'h2227: o_data_a = 16'b0000000000000000;
            14'h2228: o_data_a = 16'b1111110010100000;
            14'h2229: o_data_a = 16'b1111110001001000;
            14'h222a: o_data_a = 16'b0000000000000000;
            14'h222b: o_data_a = 16'b1111110010101000;
            14'h222c: o_data_a = 16'b1111110000010000;
            14'h222d: o_data_a = 16'b0010001001010011;
            14'h222e: o_data_a = 16'b1110001100000101;
            14'h222f: o_data_a = 16'b0000000000000000;
            14'h2230: o_data_a = 16'b1111110111001000;
            14'h2231: o_data_a = 16'b1111110010100000;
            14'h2232: o_data_a = 16'b1110111111001000;
            14'h2233: o_data_a = 16'b0000000000000001;
            14'h2234: o_data_a = 16'b1111110000100000;
            14'h2235: o_data_a = 16'b1111110000010000;
            14'h2236: o_data_a = 16'b0000000000000000;
            14'h2237: o_data_a = 16'b1111110111101000;
            14'h2238: o_data_a = 16'b1110110010100000;
            14'h2239: o_data_a = 16'b1110001100001000;
            14'h223a: o_data_a = 16'b0000000000000000;
            14'h223b: o_data_a = 16'b1111110010101000;
            14'h223c: o_data_a = 16'b1111110000010000;
            14'h223d: o_data_a = 16'b1110110010100000;
            14'h223e: o_data_a = 16'b1111000010001000;
            14'h223f: o_data_a = 16'b0000000000000000;
            14'h2240: o_data_a = 16'b1111110010101000;
            14'h2241: o_data_a = 16'b1111110000010000;
            14'h2242: o_data_a = 16'b0000000000000100;
            14'h2243: o_data_a = 16'b1110001100001000;
            14'h2244: o_data_a = 16'b0000000000000100;
            14'h2245: o_data_a = 16'b1111110000100000;
            14'h2246: o_data_a = 16'b1111110000010000;
            14'h2247: o_data_a = 16'b0000000000000000;
            14'h2248: o_data_a = 16'b1111110111101000;
            14'h2249: o_data_a = 16'b1110110010100000;
            14'h224a: o_data_a = 16'b1110001100001000;
            14'h224b: o_data_a = 16'b0000000000000000;
            14'h224c: o_data_a = 16'b1111110010101000;
            14'h224d: o_data_a = 16'b1111110000010000;
            14'h224e: o_data_a = 16'b0000000000000001;
            14'h224f: o_data_a = 16'b1111110000100000;
            14'h2250: o_data_a = 16'b1110001100001000;
            14'h2251: o_data_a = 16'b0010001000000000;
            14'h2252: o_data_a = 16'b1110101010000111;
            14'h2253: o_data_a = 16'b0000000000000001;
            14'h2254: o_data_a = 16'b1111110000100000;
            14'h2255: o_data_a = 16'b1111110000010000;
            14'h2256: o_data_a = 16'b0000000000000000;
            14'h2257: o_data_a = 16'b1111110111101000;
            14'h2258: o_data_a = 16'b1110110010100000;
            14'h2259: o_data_a = 16'b1110001100001000;
            14'h225a: o_data_a = 16'b0000000000000010;
            14'h225b: o_data_a = 16'b1111110000100000;
            14'h225c: o_data_a = 16'b1111110000010000;
            14'h225d: o_data_a = 16'b0000000000000000;
            14'h225e: o_data_a = 16'b1111110111101000;
            14'h225f: o_data_a = 16'b1110110010100000;
            14'h2260: o_data_a = 16'b1110001100001000;
            14'h2261: o_data_a = 16'b0000000000000000;
            14'h2262: o_data_a = 16'b1111110010101000;
            14'h2263: o_data_a = 16'b1111110000010000;
            14'h2264: o_data_a = 16'b1110110010100000;
            14'h2265: o_data_a = 16'b1111000010001000;
            14'h2266: o_data_a = 16'b0011111111111011;
            14'h2267: o_data_a = 16'b1110110000010000;
            14'h2268: o_data_a = 16'b0000000000000000;
            14'h2269: o_data_a = 16'b1111110111101000;
            14'h226a: o_data_a = 16'b1110110010100000;
            14'h226b: o_data_a = 16'b1110001100001000;
            14'h226c: o_data_a = 16'b0010001001110000;
            14'h226d: o_data_a = 16'b1110110000010000;
            14'h226e: o_data_a = 16'b0000000000010110;
            14'h226f: o_data_a = 16'b1110101010000111;
            14'h2270: o_data_a = 16'b0000000000000000;
            14'h2271: o_data_a = 16'b1111110010101000;
            14'h2272: o_data_a = 16'b1111110000010000;
            14'h2273: o_data_a = 16'b0010001001110111;
            14'h2274: o_data_a = 16'b1110001100000101;
            14'h2275: o_data_a = 16'b0010001010001110;
            14'h2276: o_data_a = 16'b1110101010000111;
            14'h2277: o_data_a = 16'b0000000000000110;
            14'h2278: o_data_a = 16'b1110110000010000;
            14'h2279: o_data_a = 16'b0000000000000000;
            14'h227a: o_data_a = 16'b1111110111101000;
            14'h227b: o_data_a = 16'b1110110010100000;
            14'h227c: o_data_a = 16'b1110001100001000;
            14'h227d: o_data_a = 16'b0000000000000001;
            14'h227e: o_data_a = 16'b1110110000010000;
            14'h227f: o_data_a = 16'b0000000000001101;
            14'h2280: o_data_a = 16'b1110001100001000;
            14'h2281: o_data_a = 16'b0110101011011001;
            14'h2282: o_data_a = 16'b1110110000010000;
            14'h2283: o_data_a = 16'b0000000000001110;
            14'h2284: o_data_a = 16'b1110001100001000;
            14'h2285: o_data_a = 16'b0010001010001001;
            14'h2286: o_data_a = 16'b1110110000010000;
            14'h2287: o_data_a = 16'b0000000001011111;
            14'h2288: o_data_a = 16'b1110101010000111;
            14'h2289: o_data_a = 16'b0000000000000000;
            14'h228a: o_data_a = 16'b1111110010101000;
            14'h228b: o_data_a = 16'b1111110000010000;
            14'h228c: o_data_a = 16'b0000000000000101;
            14'h228d: o_data_a = 16'b1110001100001000;
            14'h228e: o_data_a = 16'b0000000000000000;
            14'h228f: o_data_a = 16'b1111110111001000;
            14'h2290: o_data_a = 16'b1111110010100000;
            14'h2291: o_data_a = 16'b1110101010001000;
            14'h2292: o_data_a = 16'b0000000000000001;
            14'h2293: o_data_a = 16'b1111110000100000;
            14'h2294: o_data_a = 16'b1111110000010000;
            14'h2295: o_data_a = 16'b0000000000000000;
            14'h2296: o_data_a = 16'b1111110111101000;
            14'h2297: o_data_a = 16'b1110110010100000;
            14'h2298: o_data_a = 16'b1110001100001000;
            14'h2299: o_data_a = 16'b0000000000000000;
            14'h229a: o_data_a = 16'b1111110010101000;
            14'h229b: o_data_a = 16'b1111110000010000;
            14'h229c: o_data_a = 16'b1110110010100000;
            14'h229d: o_data_a = 16'b1111000010001000;
            14'h229e: o_data_a = 16'b0000000000000000;
            14'h229f: o_data_a = 16'b1111110010101000;
            14'h22a0: o_data_a = 16'b1111110000010000;
            14'h22a1: o_data_a = 16'b0000000000000100;
            14'h22a2: o_data_a = 16'b1110001100001000;
            14'h22a3: o_data_a = 16'b0000000000000100;
            14'h22a4: o_data_a = 16'b1111110000100000;
            14'h22a5: o_data_a = 16'b1111110000010000;
            14'h22a6: o_data_a = 16'b0000000000000000;
            14'h22a7: o_data_a = 16'b1111110111101000;
            14'h22a8: o_data_a = 16'b1110110010100000;
            14'h22a9: o_data_a = 16'b1110001100001000;
            14'h22aa: o_data_a = 16'b0000000000000010;
            14'h22ab: o_data_a = 16'b1111110000100000;
            14'h22ac: o_data_a = 16'b1111110000010000;
            14'h22ad: o_data_a = 16'b0000000000000000;
            14'h22ae: o_data_a = 16'b1111110111101000;
            14'h22af: o_data_a = 16'b1110110010100000;
            14'h22b0: o_data_a = 16'b1110001100001000;
            14'h22b1: o_data_a = 16'b0000000000000010;
            14'h22b2: o_data_a = 16'b1110110000010000;
            14'h22b3: o_data_a = 16'b0000000000000000;
            14'h22b4: o_data_a = 16'b1111110111101000;
            14'h22b5: o_data_a = 16'b1110110010100000;
            14'h22b6: o_data_a = 16'b1110001100001000;
            14'h22b7: o_data_a = 16'b0000000000000000;
            14'h22b8: o_data_a = 16'b1111110010101000;
            14'h22b9: o_data_a = 16'b1111110000010000;
            14'h22ba: o_data_a = 16'b1110110010100000;
            14'h22bb: o_data_a = 16'b1111000010001000;
            14'h22bc: o_data_a = 16'b0010001011000000;
            14'h22bd: o_data_a = 16'b1110110000010000;
            14'h22be: o_data_a = 16'b0000000000010110;
            14'h22bf: o_data_a = 16'b1110101010000111;
            14'h22c0: o_data_a = 16'b0000000000000000;
            14'h22c1: o_data_a = 16'b1111110010101000;
            14'h22c2: o_data_a = 16'b1111110000010000;
            14'h22c3: o_data_a = 16'b0010001011000111;
            14'h22c4: o_data_a = 16'b1110001100000101;
            14'h22c5: o_data_a = 16'b0010010001001111;
            14'h22c6: o_data_a = 16'b1110101010000111;
            14'h22c7: o_data_a = 16'b0000000000000010;
            14'h22c8: o_data_a = 16'b1111110000100000;
            14'h22c9: o_data_a = 16'b1111110000010000;
            14'h22ca: o_data_a = 16'b0000000000000000;
            14'h22cb: o_data_a = 16'b1111110111101000;
            14'h22cc: o_data_a = 16'b1110110010100000;
            14'h22cd: o_data_a = 16'b1110001100001000;
            14'h22ce: o_data_a = 16'b0000000000000010;
            14'h22cf: o_data_a = 16'b1110110000010000;
            14'h22d0: o_data_a = 16'b0000000000000000;
            14'h22d1: o_data_a = 16'b1111110111101000;
            14'h22d2: o_data_a = 16'b1110110010100000;
            14'h22d3: o_data_a = 16'b1110001100001000;
            14'h22d4: o_data_a = 16'b0000000000000000;
            14'h22d5: o_data_a = 16'b1111110010101000;
            14'h22d6: o_data_a = 16'b1111110000010000;
            14'h22d7: o_data_a = 16'b1110110010100000;
            14'h22d8: o_data_a = 16'b1111000010001000;
            14'h22d9: o_data_a = 16'b0000000000000001;
            14'h22da: o_data_a = 16'b1111110000100000;
            14'h22db: o_data_a = 16'b1111110000010000;
            14'h22dc: o_data_a = 16'b0000000000000000;
            14'h22dd: o_data_a = 16'b1111110111101000;
            14'h22de: o_data_a = 16'b1110110010100000;
            14'h22df: o_data_a = 16'b1110001100001000;
            14'h22e0: o_data_a = 16'b0000000000000000;
            14'h22e1: o_data_a = 16'b1111110010101000;
            14'h22e2: o_data_a = 16'b1111110000010000;
            14'h22e3: o_data_a = 16'b1110110010100000;
            14'h22e4: o_data_a = 16'b1111000010001000;
            14'h22e5: o_data_a = 16'b0000000000000000;
            14'h22e6: o_data_a = 16'b1111110111001000;
            14'h22e7: o_data_a = 16'b1111110010100000;
            14'h22e8: o_data_a = 16'b1110101010001000;
            14'h22e9: o_data_a = 16'b0000000000000001;
            14'h22ea: o_data_a = 16'b1111110000100000;
            14'h22eb: o_data_a = 16'b1111110000010000;
            14'h22ec: o_data_a = 16'b0000000000000000;
            14'h22ed: o_data_a = 16'b1111110111101000;
            14'h22ee: o_data_a = 16'b1110110010100000;
            14'h22ef: o_data_a = 16'b1110001100001000;
            14'h22f0: o_data_a = 16'b0000000000000000;
            14'h22f1: o_data_a = 16'b1111110010101000;
            14'h22f2: o_data_a = 16'b1111110000010000;
            14'h22f3: o_data_a = 16'b1110110010100000;
            14'h22f4: o_data_a = 16'b1111000010001000;
            14'h22f5: o_data_a = 16'b0000000000000000;
            14'h22f6: o_data_a = 16'b1111110010101000;
            14'h22f7: o_data_a = 16'b1111110000010000;
            14'h22f8: o_data_a = 16'b0000000000000100;
            14'h22f9: o_data_a = 16'b1110001100001000;
            14'h22fa: o_data_a = 16'b0000000000000100;
            14'h22fb: o_data_a = 16'b1111110000100000;
            14'h22fc: o_data_a = 16'b1111110000010000;
            14'h22fd: o_data_a = 16'b0000000000000000;
            14'h22fe: o_data_a = 16'b1111110111101000;
            14'h22ff: o_data_a = 16'b1110110010100000;
            14'h2300: o_data_a = 16'b1110001100001000;
            14'h2301: o_data_a = 16'b0000000000000010;
            14'h2302: o_data_a = 16'b1111110000100000;
            14'h2303: o_data_a = 16'b1111110000010000;
            14'h2304: o_data_a = 16'b0000000000000000;
            14'h2305: o_data_a = 16'b1111110111101000;
            14'h2306: o_data_a = 16'b1110110010100000;
            14'h2307: o_data_a = 16'b1110001100001000;
            14'h2308: o_data_a = 16'b0000000000000000;
            14'h2309: o_data_a = 16'b1111110010101000;
            14'h230a: o_data_a = 16'b1111110000010000;
            14'h230b: o_data_a = 16'b1110110010100000;
            14'h230c: o_data_a = 16'b1111000111001000;
            14'h230d: o_data_a = 16'b0000000000000010;
            14'h230e: o_data_a = 16'b1110110000010000;
            14'h230f: o_data_a = 16'b0000000000000000;
            14'h2310: o_data_a = 16'b1111110111101000;
            14'h2311: o_data_a = 16'b1110110010100000;
            14'h2312: o_data_a = 16'b1110001100001000;
            14'h2313: o_data_a = 16'b0000000000000000;
            14'h2314: o_data_a = 16'b1111110010101000;
            14'h2315: o_data_a = 16'b1111110000010000;
            14'h2316: o_data_a = 16'b1110110010100000;
            14'h2317: o_data_a = 16'b1111000111001000;
            14'h2318: o_data_a = 16'b0000000000000000;
            14'h2319: o_data_a = 16'b1111110010101000;
            14'h231a: o_data_a = 16'b1111110000010000;
            14'h231b: o_data_a = 16'b0000000000000101;
            14'h231c: o_data_a = 16'b1110001100001000;
            14'h231d: o_data_a = 16'b0000000000000000;
            14'h231e: o_data_a = 16'b1111110010101000;
            14'h231f: o_data_a = 16'b1111110000010000;
            14'h2320: o_data_a = 16'b0000000000000100;
            14'h2321: o_data_a = 16'b1110001100001000;
            14'h2322: o_data_a = 16'b0000000000000101;
            14'h2323: o_data_a = 16'b1111110000010000;
            14'h2324: o_data_a = 16'b0000000000000000;
            14'h2325: o_data_a = 16'b1111110111101000;
            14'h2326: o_data_a = 16'b1110110010100000;
            14'h2327: o_data_a = 16'b1110001100001000;
            14'h2328: o_data_a = 16'b0000000000000000;
            14'h2329: o_data_a = 16'b1111110010101000;
            14'h232a: o_data_a = 16'b1111110000010000;
            14'h232b: o_data_a = 16'b0000000000000100;
            14'h232c: o_data_a = 16'b1111110000100000;
            14'h232d: o_data_a = 16'b1110001100001000;
            14'h232e: o_data_a = 16'b0000000000000000;
            14'h232f: o_data_a = 16'b1111110111001000;
            14'h2330: o_data_a = 16'b1111110010100000;
            14'h2331: o_data_a = 16'b1110111111001000;
            14'h2332: o_data_a = 16'b0000000000000001;
            14'h2333: o_data_a = 16'b1111110000100000;
            14'h2334: o_data_a = 16'b1111110000010000;
            14'h2335: o_data_a = 16'b0000000000000000;
            14'h2336: o_data_a = 16'b1111110111101000;
            14'h2337: o_data_a = 16'b1110110010100000;
            14'h2338: o_data_a = 16'b1110001100001000;
            14'h2339: o_data_a = 16'b0000000000000000;
            14'h233a: o_data_a = 16'b1111110010101000;
            14'h233b: o_data_a = 16'b1111110000010000;
            14'h233c: o_data_a = 16'b1110110010100000;
            14'h233d: o_data_a = 16'b1111000010001000;
            14'h233e: o_data_a = 16'b0000000000000000;
            14'h233f: o_data_a = 16'b1111110010101000;
            14'h2340: o_data_a = 16'b1111110000010000;
            14'h2341: o_data_a = 16'b0000000000000100;
            14'h2342: o_data_a = 16'b1110001100001000;
            14'h2343: o_data_a = 16'b0000000000000100;
            14'h2344: o_data_a = 16'b1111110000100000;
            14'h2345: o_data_a = 16'b1111110000010000;
            14'h2346: o_data_a = 16'b0000000000000000;
            14'h2347: o_data_a = 16'b1111110111101000;
            14'h2348: o_data_a = 16'b1110110010100000;
            14'h2349: o_data_a = 16'b1110001100001000;
            14'h234a: o_data_a = 16'b0000000000000001;
            14'h234b: o_data_a = 16'b1111110000100000;
            14'h234c: o_data_a = 16'b1111110000010000;
            14'h234d: o_data_a = 16'b0000000000000000;
            14'h234e: o_data_a = 16'b1111110111101000;
            14'h234f: o_data_a = 16'b1110110010100000;
            14'h2350: o_data_a = 16'b1110001100001000;
            14'h2351: o_data_a = 16'b0000000000000010;
            14'h2352: o_data_a = 16'b1110110000010000;
            14'h2353: o_data_a = 16'b0000000000000000;
            14'h2354: o_data_a = 16'b1111110111101000;
            14'h2355: o_data_a = 16'b1110110010100000;
            14'h2356: o_data_a = 16'b1110001100001000;
            14'h2357: o_data_a = 16'b0000000000000000;
            14'h2358: o_data_a = 16'b1111110010101000;
            14'h2359: o_data_a = 16'b1111110000010000;
            14'h235a: o_data_a = 16'b1110110010100000;
            14'h235b: o_data_a = 16'b1111000010001000;
            14'h235c: o_data_a = 16'b0010001101100000;
            14'h235d: o_data_a = 16'b1110110000010000;
            14'h235e: o_data_a = 16'b0000000000000110;
            14'h235f: o_data_a = 16'b1110101010000111;
            14'h2360: o_data_a = 16'b0000000000000000;
            14'h2361: o_data_a = 16'b1111110010101000;
            14'h2362: o_data_a = 16'b1111110000010000;
            14'h2363: o_data_a = 16'b0010001101100111;
            14'h2364: o_data_a = 16'b1110001100000101;
            14'h2365: o_data_a = 16'b0010001110111011;
            14'h2366: o_data_a = 16'b1110101010000111;
            14'h2367: o_data_a = 16'b0000000000000010;
            14'h2368: o_data_a = 16'b1111110000100000;
            14'h2369: o_data_a = 16'b1111110000010000;
            14'h236a: o_data_a = 16'b0000000000000000;
            14'h236b: o_data_a = 16'b1111110111101000;
            14'h236c: o_data_a = 16'b1110110010100000;
            14'h236d: o_data_a = 16'b1110001100001000;
            14'h236e: o_data_a = 16'b0000000000000011;
            14'h236f: o_data_a = 16'b1110110000010000;
            14'h2370: o_data_a = 16'b0000000000000000;
            14'h2371: o_data_a = 16'b1111110111101000;
            14'h2372: o_data_a = 16'b1110110010100000;
            14'h2373: o_data_a = 16'b1110001100001000;
            14'h2374: o_data_a = 16'b0000000000000000;
            14'h2375: o_data_a = 16'b1111110010101000;
            14'h2376: o_data_a = 16'b1111110000010000;
            14'h2377: o_data_a = 16'b1110110010100000;
            14'h2378: o_data_a = 16'b1111000010001000;
            14'h2379: o_data_a = 16'b0000000000000001;
            14'h237a: o_data_a = 16'b1111110000100000;
            14'h237b: o_data_a = 16'b1111110000010000;
            14'h237c: o_data_a = 16'b0000000000000000;
            14'h237d: o_data_a = 16'b1111110111101000;
            14'h237e: o_data_a = 16'b1110110010100000;
            14'h237f: o_data_a = 16'b1110001100001000;
            14'h2380: o_data_a = 16'b0000000000000000;
            14'h2381: o_data_a = 16'b1111110010101000;
            14'h2382: o_data_a = 16'b1111110000010000;
            14'h2383: o_data_a = 16'b1110110010100000;
            14'h2384: o_data_a = 16'b1111000010001000;
            14'h2385: o_data_a = 16'b0000000000000001;
            14'h2386: o_data_a = 16'b1111110000100000;
            14'h2387: o_data_a = 16'b1111110000010000;
            14'h2388: o_data_a = 16'b0000000000000000;
            14'h2389: o_data_a = 16'b1111110111101000;
            14'h238a: o_data_a = 16'b1110110010100000;
            14'h238b: o_data_a = 16'b1110001100001000;
            14'h238c: o_data_a = 16'b0000000000000010;
            14'h238d: o_data_a = 16'b1111110000100000;
            14'h238e: o_data_a = 16'b1111110000010000;
            14'h238f: o_data_a = 16'b0000000000000000;
            14'h2390: o_data_a = 16'b1111110111101000;
            14'h2391: o_data_a = 16'b1110110010100000;
            14'h2392: o_data_a = 16'b1110001100001000;
            14'h2393: o_data_a = 16'b0000000000000000;
            14'h2394: o_data_a = 16'b1111110010101000;
            14'h2395: o_data_a = 16'b1111110000010000;
            14'h2396: o_data_a = 16'b1110110010100000;
            14'h2397: o_data_a = 16'b1111000010001000;
            14'h2398: o_data_a = 16'b0000000000000100;
            14'h2399: o_data_a = 16'b1110110000010000;
            14'h239a: o_data_a = 16'b0000000000000000;
            14'h239b: o_data_a = 16'b1111110111101000;
            14'h239c: o_data_a = 16'b1110110010100000;
            14'h239d: o_data_a = 16'b1110001100001000;
            14'h239e: o_data_a = 16'b0000000000000000;
            14'h239f: o_data_a = 16'b1111110010101000;
            14'h23a0: o_data_a = 16'b1111110000010000;
            14'h23a1: o_data_a = 16'b1110110010100000;
            14'h23a2: o_data_a = 16'b1111000010001000;
            14'h23a3: o_data_a = 16'b0000000000000000;
            14'h23a4: o_data_a = 16'b1111110010101000;
            14'h23a5: o_data_a = 16'b1111110000010000;
            14'h23a6: o_data_a = 16'b0000000000000101;
            14'h23a7: o_data_a = 16'b1110001100001000;
            14'h23a8: o_data_a = 16'b0000000000000000;
            14'h23a9: o_data_a = 16'b1111110010101000;
            14'h23aa: o_data_a = 16'b1111110000010000;
            14'h23ab: o_data_a = 16'b0000000000000100;
            14'h23ac: o_data_a = 16'b1110001100001000;
            14'h23ad: o_data_a = 16'b0000000000000101;
            14'h23ae: o_data_a = 16'b1111110000010000;
            14'h23af: o_data_a = 16'b0000000000000000;
            14'h23b0: o_data_a = 16'b1111110111101000;
            14'h23b1: o_data_a = 16'b1110110010100000;
            14'h23b2: o_data_a = 16'b1110001100001000;
            14'h23b3: o_data_a = 16'b0000000000000000;
            14'h23b4: o_data_a = 16'b1111110010101000;
            14'h23b5: o_data_a = 16'b1111110000010000;
            14'h23b6: o_data_a = 16'b0000000000000100;
            14'h23b7: o_data_a = 16'b1111110000100000;
            14'h23b8: o_data_a = 16'b1110001100001000;
            14'h23b9: o_data_a = 16'b0010010000001011;
            14'h23ba: o_data_a = 16'b1110101010000111;
            14'h23bb: o_data_a = 16'b0000000000000010;
            14'h23bc: o_data_a = 16'b1111110000100000;
            14'h23bd: o_data_a = 16'b1111110000010000;
            14'h23be: o_data_a = 16'b0000000000000000;
            14'h23bf: o_data_a = 16'b1111110111101000;
            14'h23c0: o_data_a = 16'b1110110010100000;
            14'h23c1: o_data_a = 16'b1110001100001000;
            14'h23c2: o_data_a = 16'b0000000000000011;
            14'h23c3: o_data_a = 16'b1110110000010000;
            14'h23c4: o_data_a = 16'b0000000000000000;
            14'h23c5: o_data_a = 16'b1111110111101000;
            14'h23c6: o_data_a = 16'b1110110010100000;
            14'h23c7: o_data_a = 16'b1110001100001000;
            14'h23c8: o_data_a = 16'b0000000000000000;
            14'h23c9: o_data_a = 16'b1111110010101000;
            14'h23ca: o_data_a = 16'b1111110000010000;
            14'h23cb: o_data_a = 16'b1110110010100000;
            14'h23cc: o_data_a = 16'b1111000010001000;
            14'h23cd: o_data_a = 16'b0000000000000001;
            14'h23ce: o_data_a = 16'b1111110000100000;
            14'h23cf: o_data_a = 16'b1111110000010000;
            14'h23d0: o_data_a = 16'b0000000000000000;
            14'h23d1: o_data_a = 16'b1111110111101000;
            14'h23d2: o_data_a = 16'b1110110010100000;
            14'h23d3: o_data_a = 16'b1110001100001000;
            14'h23d4: o_data_a = 16'b0000000000000000;
            14'h23d5: o_data_a = 16'b1111110010101000;
            14'h23d6: o_data_a = 16'b1111110000010000;
            14'h23d7: o_data_a = 16'b1110110010100000;
            14'h23d8: o_data_a = 16'b1111000010001000;
            14'h23d9: o_data_a = 16'b0000000000000000;
            14'h23da: o_data_a = 16'b1111110111001000;
            14'h23db: o_data_a = 16'b1111110010100000;
            14'h23dc: o_data_a = 16'b1110111111001000;
            14'h23dd: o_data_a = 16'b0000000000000001;
            14'h23de: o_data_a = 16'b1111110000100000;
            14'h23df: o_data_a = 16'b1111110000010000;
            14'h23e0: o_data_a = 16'b0000000000000000;
            14'h23e1: o_data_a = 16'b1111110111101000;
            14'h23e2: o_data_a = 16'b1110110010100000;
            14'h23e3: o_data_a = 16'b1110001100001000;
            14'h23e4: o_data_a = 16'b0000000000000000;
            14'h23e5: o_data_a = 16'b1111110010101000;
            14'h23e6: o_data_a = 16'b1111110000010000;
            14'h23e7: o_data_a = 16'b1110110010100000;
            14'h23e8: o_data_a = 16'b1111000010001000;
            14'h23e9: o_data_a = 16'b0000000000000000;
            14'h23ea: o_data_a = 16'b1111110010101000;
            14'h23eb: o_data_a = 16'b1111110000010000;
            14'h23ec: o_data_a = 16'b0000000000000100;
            14'h23ed: o_data_a = 16'b1110001100001000;
            14'h23ee: o_data_a = 16'b0000000000000100;
            14'h23ef: o_data_a = 16'b1111110000100000;
            14'h23f0: o_data_a = 16'b1111110000010000;
            14'h23f1: o_data_a = 16'b0000000000000000;
            14'h23f2: o_data_a = 16'b1111110111101000;
            14'h23f3: o_data_a = 16'b1110110010100000;
            14'h23f4: o_data_a = 16'b1110001100001000;
            14'h23f5: o_data_a = 16'b0000000000000000;
            14'h23f6: o_data_a = 16'b1111110010101000;
            14'h23f7: o_data_a = 16'b1111110000010000;
            14'h23f8: o_data_a = 16'b0000000000000101;
            14'h23f9: o_data_a = 16'b1110001100001000;
            14'h23fa: o_data_a = 16'b0000000000000000;
            14'h23fb: o_data_a = 16'b1111110010101000;
            14'h23fc: o_data_a = 16'b1111110000010000;
            14'h23fd: o_data_a = 16'b0000000000000100;
            14'h23fe: o_data_a = 16'b1110001100001000;
            14'h23ff: o_data_a = 16'b0000000000000101;
            14'h2400: o_data_a = 16'b1111110000010000;
            14'h2401: o_data_a = 16'b0000000000000000;
            14'h2402: o_data_a = 16'b1111110111101000;
            14'h2403: o_data_a = 16'b1110110010100000;
            14'h2404: o_data_a = 16'b1110001100001000;
            14'h2405: o_data_a = 16'b0000000000000000;
            14'h2406: o_data_a = 16'b1111110010101000;
            14'h2407: o_data_a = 16'b1111110000010000;
            14'h2408: o_data_a = 16'b0000000000000100;
            14'h2409: o_data_a = 16'b1111110000100000;
            14'h240a: o_data_a = 16'b1110001100001000;
            14'h240b: o_data_a = 16'b0000000000000000;
            14'h240c: o_data_a = 16'b1111110111001000;
            14'h240d: o_data_a = 16'b1111110010100000;
            14'h240e: o_data_a = 16'b1110111111001000;
            14'h240f: o_data_a = 16'b0000000000000001;
            14'h2410: o_data_a = 16'b1111110000100000;
            14'h2411: o_data_a = 16'b1111110000010000;
            14'h2412: o_data_a = 16'b0000000000000000;
            14'h2413: o_data_a = 16'b1111110111101000;
            14'h2414: o_data_a = 16'b1110110010100000;
            14'h2415: o_data_a = 16'b1110001100001000;
            14'h2416: o_data_a = 16'b0000000000000000;
            14'h2417: o_data_a = 16'b1111110010101000;
            14'h2418: o_data_a = 16'b1111110000010000;
            14'h2419: o_data_a = 16'b1110110010100000;
            14'h241a: o_data_a = 16'b1111000010001000;
            14'h241b: o_data_a = 16'b0000000000000001;
            14'h241c: o_data_a = 16'b1111110000100000;
            14'h241d: o_data_a = 16'b1111110000010000;
            14'h241e: o_data_a = 16'b0000000000000000;
            14'h241f: o_data_a = 16'b1111110111101000;
            14'h2420: o_data_a = 16'b1110110010100000;
            14'h2421: o_data_a = 16'b1110001100001000;
            14'h2422: o_data_a = 16'b0000000000000010;
            14'h2423: o_data_a = 16'b1111110000100000;
            14'h2424: o_data_a = 16'b1111110000010000;
            14'h2425: o_data_a = 16'b0000000000000000;
            14'h2426: o_data_a = 16'b1111110111101000;
            14'h2427: o_data_a = 16'b1110110010100000;
            14'h2428: o_data_a = 16'b1110001100001000;
            14'h2429: o_data_a = 16'b0000000000000000;
            14'h242a: o_data_a = 16'b1111110010101000;
            14'h242b: o_data_a = 16'b1111110000010000;
            14'h242c: o_data_a = 16'b1110110010100000;
            14'h242d: o_data_a = 16'b1111000010001000;
            14'h242e: o_data_a = 16'b0000000000000010;
            14'h242f: o_data_a = 16'b1110110000010000;
            14'h2430: o_data_a = 16'b0000000000000000;
            14'h2431: o_data_a = 16'b1111110111101000;
            14'h2432: o_data_a = 16'b1110110010100000;
            14'h2433: o_data_a = 16'b1110001100001000;
            14'h2434: o_data_a = 16'b0000000000000000;
            14'h2435: o_data_a = 16'b1111110010101000;
            14'h2436: o_data_a = 16'b1111110000010000;
            14'h2437: o_data_a = 16'b1110110010100000;
            14'h2438: o_data_a = 16'b1111000010001000;
            14'h2439: o_data_a = 16'b0000000000000000;
            14'h243a: o_data_a = 16'b1111110010101000;
            14'h243b: o_data_a = 16'b1111110000010000;
            14'h243c: o_data_a = 16'b0000000000000101;
            14'h243d: o_data_a = 16'b1110001100001000;
            14'h243e: o_data_a = 16'b0000000000000000;
            14'h243f: o_data_a = 16'b1111110010101000;
            14'h2440: o_data_a = 16'b1111110000010000;
            14'h2441: o_data_a = 16'b0000000000000100;
            14'h2442: o_data_a = 16'b1110001100001000;
            14'h2443: o_data_a = 16'b0000000000000101;
            14'h2444: o_data_a = 16'b1111110000010000;
            14'h2445: o_data_a = 16'b0000000000000000;
            14'h2446: o_data_a = 16'b1111110111101000;
            14'h2447: o_data_a = 16'b1110110010100000;
            14'h2448: o_data_a = 16'b1110001100001000;
            14'h2449: o_data_a = 16'b0000000000000000;
            14'h244a: o_data_a = 16'b1111110010101000;
            14'h244b: o_data_a = 16'b1111110000010000;
            14'h244c: o_data_a = 16'b0000000000000100;
            14'h244d: o_data_a = 16'b1111110000100000;
            14'h244e: o_data_a = 16'b1110001100001000;
            14'h244f: o_data_a = 16'b0000000000000000;
            14'h2450: o_data_a = 16'b1111110111001000;
            14'h2451: o_data_a = 16'b1111110010100000;
            14'h2452: o_data_a = 16'b1110101010001000;
            14'h2453: o_data_a = 16'b0000000000000001;
            14'h2454: o_data_a = 16'b1111110000100000;
            14'h2455: o_data_a = 16'b1111110000010000;
            14'h2456: o_data_a = 16'b0000000000000000;
            14'h2457: o_data_a = 16'b1111110111101000;
            14'h2458: o_data_a = 16'b1110110010100000;
            14'h2459: o_data_a = 16'b1110001100001000;
            14'h245a: o_data_a = 16'b0000000000000000;
            14'h245b: o_data_a = 16'b1111110010101000;
            14'h245c: o_data_a = 16'b1111110000010000;
            14'h245d: o_data_a = 16'b1110110010100000;
            14'h245e: o_data_a = 16'b1111000010001000;
            14'h245f: o_data_a = 16'b0000000000000000;
            14'h2460: o_data_a = 16'b1111110111001000;
            14'h2461: o_data_a = 16'b1111110010100000;
            14'h2462: o_data_a = 16'b1110101010001000;
            14'h2463: o_data_a = 16'b0000000000000000;
            14'h2464: o_data_a = 16'b1111110010101000;
            14'h2465: o_data_a = 16'b1111110000010000;
            14'h2466: o_data_a = 16'b0000000000000101;
            14'h2467: o_data_a = 16'b1110001100001000;
            14'h2468: o_data_a = 16'b0000000000000000;
            14'h2469: o_data_a = 16'b1111110010101000;
            14'h246a: o_data_a = 16'b1111110000010000;
            14'h246b: o_data_a = 16'b0000000000000100;
            14'h246c: o_data_a = 16'b1110001100001000;
            14'h246d: o_data_a = 16'b0000000000000101;
            14'h246e: o_data_a = 16'b1111110000010000;
            14'h246f: o_data_a = 16'b0000000000000000;
            14'h2470: o_data_a = 16'b1111110111101000;
            14'h2471: o_data_a = 16'b1110110010100000;
            14'h2472: o_data_a = 16'b1110001100001000;
            14'h2473: o_data_a = 16'b0000000000000000;
            14'h2474: o_data_a = 16'b1111110010101000;
            14'h2475: o_data_a = 16'b1111110000010000;
            14'h2476: o_data_a = 16'b0000000000000100;
            14'h2477: o_data_a = 16'b1111110000100000;
            14'h2478: o_data_a = 16'b1110001100001000;
            14'h2479: o_data_a = 16'b0000000000000001;
            14'h247a: o_data_a = 16'b1111110000100000;
            14'h247b: o_data_a = 16'b1111110000010000;
            14'h247c: o_data_a = 16'b0000000000000000;
            14'h247d: o_data_a = 16'b1111110111101000;
            14'h247e: o_data_a = 16'b1110110010100000;
            14'h247f: o_data_a = 16'b1110001100001000;
            14'h2480: o_data_a = 16'b0000000000000010;
            14'h2481: o_data_a = 16'b1110110000010000;
            14'h2482: o_data_a = 16'b0000000000000000;
            14'h2483: o_data_a = 16'b1111110111101000;
            14'h2484: o_data_a = 16'b1110110010100000;
            14'h2485: o_data_a = 16'b1110001100001000;
            14'h2486: o_data_a = 16'b0000000000000000;
            14'h2487: o_data_a = 16'b1111110010101000;
            14'h2488: o_data_a = 16'b1111110000010000;
            14'h2489: o_data_a = 16'b1110110010100000;
            14'h248a: o_data_a = 16'b1111000010001000;
            14'h248b: o_data_a = 16'b0000000000110110;
            14'h248c: o_data_a = 16'b1110101010000111;
            14'h248d: o_data_a = 16'b0000000000000000;
            14'h248e: o_data_a = 16'b1111110000100000;
            14'h248f: o_data_a = 16'b1110101010001000;
            14'h2490: o_data_a = 16'b1110110111110000;
            14'h2491: o_data_a = 16'b1110101010001000;
            14'h2492: o_data_a = 16'b0000000000000000;
            14'h2493: o_data_a = 16'b1110011111001000;
            14'h2494: o_data_a = 16'b0000000000000010;
            14'h2495: o_data_a = 16'b1111110000100000;
            14'h2496: o_data_a = 16'b1111110000010000;
            14'h2497: o_data_a = 16'b0000000000000000;
            14'h2498: o_data_a = 16'b1111110111101000;
            14'h2499: o_data_a = 16'b1110110010100000;
            14'h249a: o_data_a = 16'b1110001100001000;
            14'h249b: o_data_a = 16'b0000000000000010;
            14'h249c: o_data_a = 16'b1110110000010000;
            14'h249d: o_data_a = 16'b0000000000000000;
            14'h249e: o_data_a = 16'b1111110111101000;
            14'h249f: o_data_a = 16'b1110110010100000;
            14'h24a0: o_data_a = 16'b1110001100001000;
            14'h24a1: o_data_a = 16'b0000000000000000;
            14'h24a2: o_data_a = 16'b1111110010101000;
            14'h24a3: o_data_a = 16'b1111110000010000;
            14'h24a4: o_data_a = 16'b1110110010100000;
            14'h24a5: o_data_a = 16'b1111000111001000;
            14'h24a6: o_data_a = 16'b0000000000000000;
            14'h24a7: o_data_a = 16'b1111110010101000;
            14'h24a8: o_data_a = 16'b1111110000010000;
            14'h24a9: o_data_a = 16'b0000000000000001;
            14'h24aa: o_data_a = 16'b1111110000100000;
            14'h24ab: o_data_a = 16'b1110001100001000;
            14'h24ac: o_data_a = 16'b0000000000000000;
            14'h24ad: o_data_a = 16'b1111110111001000;
            14'h24ae: o_data_a = 16'b1111110010100000;
            14'h24af: o_data_a = 16'b1110111111001000;
            14'h24b0: o_data_a = 16'b0000000000000001;
            14'h24b1: o_data_a = 16'b1111110000100000;
            14'h24b2: o_data_a = 16'b1111110000010000;
            14'h24b3: o_data_a = 16'b0000000000000000;
            14'h24b4: o_data_a = 16'b1111110111101000;
            14'h24b5: o_data_a = 16'b1110110010100000;
            14'h24b6: o_data_a = 16'b1110001100001000;
            14'h24b7: o_data_a = 16'b0000000000000000;
            14'h24b8: o_data_a = 16'b1111110010101000;
            14'h24b9: o_data_a = 16'b1111110000010000;
            14'h24ba: o_data_a = 16'b1110110010100000;
            14'h24bb: o_data_a = 16'b1111000010001000;
            14'h24bc: o_data_a = 16'b0000000000000000;
            14'h24bd: o_data_a = 16'b1111110010101000;
            14'h24be: o_data_a = 16'b1111110000010000;
            14'h24bf: o_data_a = 16'b0000000000000100;
            14'h24c0: o_data_a = 16'b1110001100001000;
            14'h24c1: o_data_a = 16'b0000000000000100;
            14'h24c2: o_data_a = 16'b1111110000100000;
            14'h24c3: o_data_a = 16'b1111110000010000;
            14'h24c4: o_data_a = 16'b0000000000000000;
            14'h24c5: o_data_a = 16'b1111110111101000;
            14'h24c6: o_data_a = 16'b1110110010100000;
            14'h24c7: o_data_a = 16'b1110001100001000;
            14'h24c8: o_data_a = 16'b0000000000000000;
            14'h24c9: o_data_a = 16'b1111110010101000;
            14'h24ca: o_data_a = 16'b1111110000010000;
            14'h24cb: o_data_a = 16'b0000000000000001;
            14'h24cc: o_data_a = 16'b1111110111100000;
            14'h24cd: o_data_a = 16'b1110001100001000;
            14'h24ce: o_data_a = 16'b0000000000000000;
            14'h24cf: o_data_a = 16'b1111110111001000;
            14'h24d0: o_data_a = 16'b1111110010100000;
            14'h24d1: o_data_a = 16'b1110101010001000;
            14'h24d2: o_data_a = 16'b0000000000000001;
            14'h24d3: o_data_a = 16'b1111110111100000;
            14'h24d4: o_data_a = 16'b1111110000010000;
            14'h24d5: o_data_a = 16'b0000000000000000;
            14'h24d6: o_data_a = 16'b1111110111101000;
            14'h24d7: o_data_a = 16'b1110110010100000;
            14'h24d8: o_data_a = 16'b1110001100001000;
            14'h24d9: o_data_a = 16'b0000000000000000;
            14'h24da: o_data_a = 16'b1111110010101000;
            14'h24db: o_data_a = 16'b1111110000010000;
            14'h24dc: o_data_a = 16'b1110110010100000;
            14'h24dd: o_data_a = 16'b1111000010001000;
            14'h24de: o_data_a = 16'b0000000000000000;
            14'h24df: o_data_a = 16'b1111110010101000;
            14'h24e0: o_data_a = 16'b1111110000010000;
            14'h24e1: o_data_a = 16'b0000000000000100;
            14'h24e2: o_data_a = 16'b1110001100001000;
            14'h24e3: o_data_a = 16'b0000000000000100;
            14'h24e4: o_data_a = 16'b1111110000100000;
            14'h24e5: o_data_a = 16'b1111110000010000;
            14'h24e6: o_data_a = 16'b0000000000000000;
            14'h24e7: o_data_a = 16'b1111110111101000;
            14'h24e8: o_data_a = 16'b1110110010100000;
            14'h24e9: o_data_a = 16'b1110001100001000;
            14'h24ea: o_data_a = 16'b0000000000000000;
            14'h24eb: o_data_a = 16'b1111110111001000;
            14'h24ec: o_data_a = 16'b1111110010100000;
            14'h24ed: o_data_a = 16'b1110101010001000;
            14'h24ee: o_data_a = 16'b0010010011110010;
            14'h24ef: o_data_a = 16'b1110110000010000;
            14'h24f0: o_data_a = 16'b0000000000000110;
            14'h24f1: o_data_a = 16'b1110101010000111;
            14'h24f2: o_data_a = 16'b0000000000000000;
            14'h24f3: o_data_a = 16'b1111110010101000;
            14'h24f4: o_data_a = 16'b1111110000010000;
            14'h24f5: o_data_a = 16'b0010010011111001;
            14'h24f6: o_data_a = 16'b1110001100000101;
            14'h24f7: o_data_a = 16'b0010010101010100;
            14'h24f8: o_data_a = 16'b1110101010000111;
            14'h24f9: o_data_a = 16'b0000000000000000;
            14'h24fa: o_data_a = 16'b1111110111001000;
            14'h24fb: o_data_a = 16'b1111110010100000;
            14'h24fc: o_data_a = 16'b1110101010001000;
            14'h24fd: o_data_a = 16'b0000000000000001;
            14'h24fe: o_data_a = 16'b1111110000100000;
            14'h24ff: o_data_a = 16'b1111110000010000;
            14'h2500: o_data_a = 16'b0000000000000000;
            14'h2501: o_data_a = 16'b1111110111101000;
            14'h2502: o_data_a = 16'b1110110010100000;
            14'h2503: o_data_a = 16'b1110001100001000;
            14'h2504: o_data_a = 16'b0000000000000000;
            14'h2505: o_data_a = 16'b1111110010101000;
            14'h2506: o_data_a = 16'b1111110000010000;
            14'h2507: o_data_a = 16'b1110110010100000;
            14'h2508: o_data_a = 16'b1111000010001000;
            14'h2509: o_data_a = 16'b0000000000000000;
            14'h250a: o_data_a = 16'b1111110111001000;
            14'h250b: o_data_a = 16'b1111110010100000;
            14'h250c: o_data_a = 16'b1110111111001000;
            14'h250d: o_data_a = 16'b0000000000000001;
            14'h250e: o_data_a = 16'b1111110000100000;
            14'h250f: o_data_a = 16'b1111110000010000;
            14'h2510: o_data_a = 16'b0000000000000000;
            14'h2511: o_data_a = 16'b1111110111101000;
            14'h2512: o_data_a = 16'b1110110010100000;
            14'h2513: o_data_a = 16'b1110001100001000;
            14'h2514: o_data_a = 16'b0000000000000000;
            14'h2515: o_data_a = 16'b1111110010101000;
            14'h2516: o_data_a = 16'b1111110000010000;
            14'h2517: o_data_a = 16'b1110110010100000;
            14'h2518: o_data_a = 16'b1111000010001000;
            14'h2519: o_data_a = 16'b0000000000000000;
            14'h251a: o_data_a = 16'b1111110010101000;
            14'h251b: o_data_a = 16'b1111110000010000;
            14'h251c: o_data_a = 16'b0000000000000100;
            14'h251d: o_data_a = 16'b1110001100001000;
            14'h251e: o_data_a = 16'b0000000000000100;
            14'h251f: o_data_a = 16'b1111110000100000;
            14'h2520: o_data_a = 16'b1111110000010000;
            14'h2521: o_data_a = 16'b0000000000000000;
            14'h2522: o_data_a = 16'b1111110111101000;
            14'h2523: o_data_a = 16'b1110110010100000;
            14'h2524: o_data_a = 16'b1110001100001000;
            14'h2525: o_data_a = 16'b0000000000000001;
            14'h2526: o_data_a = 16'b1111110000100000;
            14'h2527: o_data_a = 16'b1111110000010000;
            14'h2528: o_data_a = 16'b0000000000000000;
            14'h2529: o_data_a = 16'b1111110111101000;
            14'h252a: o_data_a = 16'b1110110010100000;
            14'h252b: o_data_a = 16'b1110001100001000;
            14'h252c: o_data_a = 16'b0000000000000000;
            14'h252d: o_data_a = 16'b1111110010101000;
            14'h252e: o_data_a = 16'b1111110000010000;
            14'h252f: o_data_a = 16'b1110110010100000;
            14'h2530: o_data_a = 16'b1111000111001000;
            14'h2531: o_data_a = 16'b0000000000000010;
            14'h2532: o_data_a = 16'b1110110000010000;
            14'h2533: o_data_a = 16'b0000000000000000;
            14'h2534: o_data_a = 16'b1111110111101000;
            14'h2535: o_data_a = 16'b1110110010100000;
            14'h2536: o_data_a = 16'b1110001100001000;
            14'h2537: o_data_a = 16'b0000000000000000;
            14'h2538: o_data_a = 16'b1111110010101000;
            14'h2539: o_data_a = 16'b1111110000010000;
            14'h253a: o_data_a = 16'b1110110010100000;
            14'h253b: o_data_a = 16'b1111000111001000;
            14'h253c: o_data_a = 16'b0000000000000000;
            14'h253d: o_data_a = 16'b1111110010101000;
            14'h253e: o_data_a = 16'b1111110000010000;
            14'h253f: o_data_a = 16'b0000000000000101;
            14'h2540: o_data_a = 16'b1110001100001000;
            14'h2541: o_data_a = 16'b0000000000000000;
            14'h2542: o_data_a = 16'b1111110010101000;
            14'h2543: o_data_a = 16'b1111110000010000;
            14'h2544: o_data_a = 16'b0000000000000100;
            14'h2545: o_data_a = 16'b1110001100001000;
            14'h2546: o_data_a = 16'b0000000000000101;
            14'h2547: o_data_a = 16'b1111110000010000;
            14'h2548: o_data_a = 16'b0000000000000000;
            14'h2549: o_data_a = 16'b1111110111101000;
            14'h254a: o_data_a = 16'b1110110010100000;
            14'h254b: o_data_a = 16'b1110001100001000;
            14'h254c: o_data_a = 16'b0000000000000000;
            14'h254d: o_data_a = 16'b1111110010101000;
            14'h254e: o_data_a = 16'b1111110000010000;
            14'h254f: o_data_a = 16'b0000000000000100;
            14'h2550: o_data_a = 16'b1111110000100000;
            14'h2551: o_data_a = 16'b1110001100001000;
            14'h2552: o_data_a = 16'b0010011001111000;
            14'h2553: o_data_a = 16'b1110101010000111;
            14'h2554: o_data_a = 16'b0000000000000000;
            14'h2555: o_data_a = 16'b1111110111001000;
            14'h2556: o_data_a = 16'b1111110010100000;
            14'h2557: o_data_a = 16'b1110101010001000;
            14'h2558: o_data_a = 16'b0000000000000001;
            14'h2559: o_data_a = 16'b1111110000100000;
            14'h255a: o_data_a = 16'b1111110000010000;
            14'h255b: o_data_a = 16'b0000000000000000;
            14'h255c: o_data_a = 16'b1111110111101000;
            14'h255d: o_data_a = 16'b1110110010100000;
            14'h255e: o_data_a = 16'b1110001100001000;
            14'h255f: o_data_a = 16'b0000000000000000;
            14'h2560: o_data_a = 16'b1111110010101000;
            14'h2561: o_data_a = 16'b1111110000010000;
            14'h2562: o_data_a = 16'b1110110010100000;
            14'h2563: o_data_a = 16'b1111000010001000;
            14'h2564: o_data_a = 16'b0000000000000000;
            14'h2565: o_data_a = 16'b1111110111001000;
            14'h2566: o_data_a = 16'b1111110010100000;
            14'h2567: o_data_a = 16'b1110111111001000;
            14'h2568: o_data_a = 16'b0000000000000001;
            14'h2569: o_data_a = 16'b1111110000100000;
            14'h256a: o_data_a = 16'b1111110000010000;
            14'h256b: o_data_a = 16'b0000000000000000;
            14'h256c: o_data_a = 16'b1111110111101000;
            14'h256d: o_data_a = 16'b1110110010100000;
            14'h256e: o_data_a = 16'b1110001100001000;
            14'h256f: o_data_a = 16'b0000000000000000;
            14'h2570: o_data_a = 16'b1111110010101000;
            14'h2571: o_data_a = 16'b1111110000010000;
            14'h2572: o_data_a = 16'b1110110010100000;
            14'h2573: o_data_a = 16'b1111000010001000;
            14'h2574: o_data_a = 16'b0000000000000000;
            14'h2575: o_data_a = 16'b1111110010101000;
            14'h2576: o_data_a = 16'b1111110000010000;
            14'h2577: o_data_a = 16'b0000000000000100;
            14'h2578: o_data_a = 16'b1110001100001000;
            14'h2579: o_data_a = 16'b0000000000000100;
            14'h257a: o_data_a = 16'b1111110000100000;
            14'h257b: o_data_a = 16'b1111110000010000;
            14'h257c: o_data_a = 16'b0000000000000000;
            14'h257d: o_data_a = 16'b1111110111101000;
            14'h257e: o_data_a = 16'b1110110010100000;
            14'h257f: o_data_a = 16'b1110001100001000;
            14'h2580: o_data_a = 16'b0000000000000001;
            14'h2581: o_data_a = 16'b1111110000100000;
            14'h2582: o_data_a = 16'b1111110000010000;
            14'h2583: o_data_a = 16'b0000000000000000;
            14'h2584: o_data_a = 16'b1111110111101000;
            14'h2585: o_data_a = 16'b1110110010100000;
            14'h2586: o_data_a = 16'b1110001100001000;
            14'h2587: o_data_a = 16'b0000000000000000;
            14'h2588: o_data_a = 16'b1111110010101000;
            14'h2589: o_data_a = 16'b1111110000010000;
            14'h258a: o_data_a = 16'b1110110010100000;
            14'h258b: o_data_a = 16'b1111000111001000;
            14'h258c: o_data_a = 16'b0000000000000000;
            14'h258d: o_data_a = 16'b1111110111001000;
            14'h258e: o_data_a = 16'b1111110010100000;
            14'h258f: o_data_a = 16'b1110101010001000;
            14'h2590: o_data_a = 16'b0000000000000001;
            14'h2591: o_data_a = 16'b1111110111100000;
            14'h2592: o_data_a = 16'b1111110000010000;
            14'h2593: o_data_a = 16'b0000000000000000;
            14'h2594: o_data_a = 16'b1111110111101000;
            14'h2595: o_data_a = 16'b1110110010100000;
            14'h2596: o_data_a = 16'b1110001100001000;
            14'h2597: o_data_a = 16'b0000000000000000;
            14'h2598: o_data_a = 16'b1111110010101000;
            14'h2599: o_data_a = 16'b1111110000010000;
            14'h259a: o_data_a = 16'b1110110010100000;
            14'h259b: o_data_a = 16'b1111000010001000;
            14'h259c: o_data_a = 16'b0000000000000000;
            14'h259d: o_data_a = 16'b1111110010101000;
            14'h259e: o_data_a = 16'b1111110000010000;
            14'h259f: o_data_a = 16'b0000000000000100;
            14'h25a0: o_data_a = 16'b1110001100001000;
            14'h25a1: o_data_a = 16'b0000000000000100;
            14'h25a2: o_data_a = 16'b1111110000100000;
            14'h25a3: o_data_a = 16'b1111110000010000;
            14'h25a4: o_data_a = 16'b0000000000000000;
            14'h25a5: o_data_a = 16'b1111110111101000;
            14'h25a6: o_data_a = 16'b1110110010100000;
            14'h25a7: o_data_a = 16'b1110001100001000;
            14'h25a8: o_data_a = 16'b0000000000000000;
            14'h25a9: o_data_a = 16'b1111110010101000;
            14'h25aa: o_data_a = 16'b1111110000010000;
            14'h25ab: o_data_a = 16'b1110110010100000;
            14'h25ac: o_data_a = 16'b1111000010001000;
            14'h25ad: o_data_a = 16'b0000000000000000;
            14'h25ae: o_data_a = 16'b1111110010101000;
            14'h25af: o_data_a = 16'b1111110000010000;
            14'h25b0: o_data_a = 16'b0000000000000101;
            14'h25b1: o_data_a = 16'b1110001100001000;
            14'h25b2: o_data_a = 16'b0000000000000000;
            14'h25b3: o_data_a = 16'b1111110010101000;
            14'h25b4: o_data_a = 16'b1111110000010000;
            14'h25b5: o_data_a = 16'b0000000000000100;
            14'h25b6: o_data_a = 16'b1110001100001000;
            14'h25b7: o_data_a = 16'b0000000000000101;
            14'h25b8: o_data_a = 16'b1111110000010000;
            14'h25b9: o_data_a = 16'b0000000000000000;
            14'h25ba: o_data_a = 16'b1111110111101000;
            14'h25bb: o_data_a = 16'b1110110010100000;
            14'h25bc: o_data_a = 16'b1110001100001000;
            14'h25bd: o_data_a = 16'b0000000000000000;
            14'h25be: o_data_a = 16'b1111110010101000;
            14'h25bf: o_data_a = 16'b1111110000010000;
            14'h25c0: o_data_a = 16'b0000000000000100;
            14'h25c1: o_data_a = 16'b1111110000100000;
            14'h25c2: o_data_a = 16'b1110001100001000;
            14'h25c3: o_data_a = 16'b0000000000000000;
            14'h25c4: o_data_a = 16'b1111110111001000;
            14'h25c5: o_data_a = 16'b1111110010100000;
            14'h25c6: o_data_a = 16'b1110111111001000;
            14'h25c7: o_data_a = 16'b0000000000000001;
            14'h25c8: o_data_a = 16'b1111110111100000;
            14'h25c9: o_data_a = 16'b1111110000010000;
            14'h25ca: o_data_a = 16'b0000000000000000;
            14'h25cb: o_data_a = 16'b1111110111101000;
            14'h25cc: o_data_a = 16'b1110110010100000;
            14'h25cd: o_data_a = 16'b1110001100001000;
            14'h25ce: o_data_a = 16'b0000000000000000;
            14'h25cf: o_data_a = 16'b1111110010101000;
            14'h25d0: o_data_a = 16'b1111110000010000;
            14'h25d1: o_data_a = 16'b1110110010100000;
            14'h25d2: o_data_a = 16'b1111000010001000;
            14'h25d3: o_data_a = 16'b0000000000000000;
            14'h25d4: o_data_a = 16'b1111110010101000;
            14'h25d5: o_data_a = 16'b1111110000010000;
            14'h25d6: o_data_a = 16'b0000000000000100;
            14'h25d7: o_data_a = 16'b1110001100001000;
            14'h25d8: o_data_a = 16'b0000000000000100;
            14'h25d9: o_data_a = 16'b1111110000100000;
            14'h25da: o_data_a = 16'b1111110000010000;
            14'h25db: o_data_a = 16'b0000000000000000;
            14'h25dc: o_data_a = 16'b1111110111101000;
            14'h25dd: o_data_a = 16'b1110110010100000;
            14'h25de: o_data_a = 16'b1110001100001000;
            14'h25df: o_data_a = 16'b0000000000000001;
            14'h25e0: o_data_a = 16'b1111110111100000;
            14'h25e1: o_data_a = 16'b1111110000010000;
            14'h25e2: o_data_a = 16'b0000000000000000;
            14'h25e3: o_data_a = 16'b1111110111101000;
            14'h25e4: o_data_a = 16'b1110110010100000;
            14'h25e5: o_data_a = 16'b1110001100001000;
            14'h25e6: o_data_a = 16'b0000000000000010;
            14'h25e7: o_data_a = 16'b1110110000010000;
            14'h25e8: o_data_a = 16'b0000000000000000;
            14'h25e9: o_data_a = 16'b1111110111101000;
            14'h25ea: o_data_a = 16'b1110110010100000;
            14'h25eb: o_data_a = 16'b1110001100001000;
            14'h25ec: o_data_a = 16'b0000000000000000;
            14'h25ed: o_data_a = 16'b1111110010101000;
            14'h25ee: o_data_a = 16'b1111110000010000;
            14'h25ef: o_data_a = 16'b1110110010100000;
            14'h25f0: o_data_a = 16'b1111000010001000;
            14'h25f1: o_data_a = 16'b0010010111110101;
            14'h25f2: o_data_a = 16'b1110110000010000;
            14'h25f3: o_data_a = 16'b0000000000000110;
            14'h25f4: o_data_a = 16'b1110101010000111;
            14'h25f5: o_data_a = 16'b0000000000000000;
            14'h25f6: o_data_a = 16'b1111110010101000;
            14'h25f7: o_data_a = 16'b1111110000010000;
            14'h25f8: o_data_a = 16'b0010010111111100;
            14'h25f9: o_data_a = 16'b1110001100000101;
            14'h25fa: o_data_a = 16'b0010011000110110;
            14'h25fb: o_data_a = 16'b1110101010000111;
            14'h25fc: o_data_a = 16'b0000000000000000;
            14'h25fd: o_data_a = 16'b1111110111001000;
            14'h25fe: o_data_a = 16'b1111110010100000;
            14'h25ff: o_data_a = 16'b1110111111001000;
            14'h2600: o_data_a = 16'b0000000000000001;
            14'h2601: o_data_a = 16'b1111110000100000;
            14'h2602: o_data_a = 16'b1111110000010000;
            14'h2603: o_data_a = 16'b0000000000000000;
            14'h2604: o_data_a = 16'b1111110111101000;
            14'h2605: o_data_a = 16'b1110110010100000;
            14'h2606: o_data_a = 16'b1110001100001000;
            14'h2607: o_data_a = 16'b0000000000000000;
            14'h2608: o_data_a = 16'b1111110010101000;
            14'h2609: o_data_a = 16'b1111110000010000;
            14'h260a: o_data_a = 16'b1110110010100000;
            14'h260b: o_data_a = 16'b1111000010001000;
            14'h260c: o_data_a = 16'b0000000000000001;
            14'h260d: o_data_a = 16'b1111110000100000;
            14'h260e: o_data_a = 16'b1111110000010000;
            14'h260f: o_data_a = 16'b0000000000000000;
            14'h2610: o_data_a = 16'b1111110111101000;
            14'h2611: o_data_a = 16'b1110110010100000;
            14'h2612: o_data_a = 16'b1110001100001000;
            14'h2613: o_data_a = 16'b0000000000000010;
            14'h2614: o_data_a = 16'b1110110000010000;
            14'h2615: o_data_a = 16'b0000000000000000;
            14'h2616: o_data_a = 16'b1111110111101000;
            14'h2617: o_data_a = 16'b1110110010100000;
            14'h2618: o_data_a = 16'b1110001100001000;
            14'h2619: o_data_a = 16'b0000000000000000;
            14'h261a: o_data_a = 16'b1111110010101000;
            14'h261b: o_data_a = 16'b1111110000010000;
            14'h261c: o_data_a = 16'b1110110010100000;
            14'h261d: o_data_a = 16'b1111000010001000;
            14'h261e: o_data_a = 16'b0000000000000000;
            14'h261f: o_data_a = 16'b1111110010101000;
            14'h2620: o_data_a = 16'b1111110000010000;
            14'h2621: o_data_a = 16'b0000000000000101;
            14'h2622: o_data_a = 16'b1110001100001000;
            14'h2623: o_data_a = 16'b0000000000000000;
            14'h2624: o_data_a = 16'b1111110010101000;
            14'h2625: o_data_a = 16'b1111110000010000;
            14'h2626: o_data_a = 16'b0000000000000100;
            14'h2627: o_data_a = 16'b1110001100001000;
            14'h2628: o_data_a = 16'b0000000000000101;
            14'h2629: o_data_a = 16'b1111110000010000;
            14'h262a: o_data_a = 16'b0000000000000000;
            14'h262b: o_data_a = 16'b1111110111101000;
            14'h262c: o_data_a = 16'b1110110010100000;
            14'h262d: o_data_a = 16'b1110001100001000;
            14'h262e: o_data_a = 16'b0000000000000000;
            14'h262f: o_data_a = 16'b1111110010101000;
            14'h2630: o_data_a = 16'b1111110000010000;
            14'h2631: o_data_a = 16'b0000000000000100;
            14'h2632: o_data_a = 16'b1111110000100000;
            14'h2633: o_data_a = 16'b1110001100001000;
            14'h2634: o_data_a = 16'b0010011001111000;
            14'h2635: o_data_a = 16'b1110101010000111;
            14'h2636: o_data_a = 16'b0000000000000000;
            14'h2637: o_data_a = 16'b1111110111001000;
            14'h2638: o_data_a = 16'b1111110010100000;
            14'h2639: o_data_a = 16'b1110111111001000;
            14'h263a: o_data_a = 16'b0000000000000001;
            14'h263b: o_data_a = 16'b1111110000100000;
            14'h263c: o_data_a = 16'b1111110000010000;
            14'h263d: o_data_a = 16'b0000000000000000;
            14'h263e: o_data_a = 16'b1111110111101000;
            14'h263f: o_data_a = 16'b1110110010100000;
            14'h2640: o_data_a = 16'b1110001100001000;
            14'h2641: o_data_a = 16'b0000000000000000;
            14'h2642: o_data_a = 16'b1111110010101000;
            14'h2643: o_data_a = 16'b1111110000010000;
            14'h2644: o_data_a = 16'b1110110010100000;
            14'h2645: o_data_a = 16'b1111000010001000;
            14'h2646: o_data_a = 16'b0000000000000000;
            14'h2647: o_data_a = 16'b1111110111001000;
            14'h2648: o_data_a = 16'b1111110010100000;
            14'h2649: o_data_a = 16'b1110111111001000;
            14'h264a: o_data_a = 16'b0000000000000001;
            14'h264b: o_data_a = 16'b1111110111100000;
            14'h264c: o_data_a = 16'b1111110000010000;
            14'h264d: o_data_a = 16'b0000000000000000;
            14'h264e: o_data_a = 16'b1111110111101000;
            14'h264f: o_data_a = 16'b1110110010100000;
            14'h2650: o_data_a = 16'b1110001100001000;
            14'h2651: o_data_a = 16'b0000000000000000;
            14'h2652: o_data_a = 16'b1111110010101000;
            14'h2653: o_data_a = 16'b1111110000010000;
            14'h2654: o_data_a = 16'b1110110010100000;
            14'h2655: o_data_a = 16'b1111000010001000;
            14'h2656: o_data_a = 16'b0000000000000000;
            14'h2657: o_data_a = 16'b1111110010101000;
            14'h2658: o_data_a = 16'b1111110000010000;
            14'h2659: o_data_a = 16'b0000000000000100;
            14'h265a: o_data_a = 16'b1110001100001000;
            14'h265b: o_data_a = 16'b0000000000000100;
            14'h265c: o_data_a = 16'b1111110000100000;
            14'h265d: o_data_a = 16'b1111110000010000;
            14'h265e: o_data_a = 16'b0000000000000000;
            14'h265f: o_data_a = 16'b1111110111101000;
            14'h2660: o_data_a = 16'b1110110010100000;
            14'h2661: o_data_a = 16'b1110001100001000;
            14'h2662: o_data_a = 16'b0000000000000000;
            14'h2663: o_data_a = 16'b1111110010101000;
            14'h2664: o_data_a = 16'b1111110000010000;
            14'h2665: o_data_a = 16'b0000000000000101;
            14'h2666: o_data_a = 16'b1110001100001000;
            14'h2667: o_data_a = 16'b0000000000000000;
            14'h2668: o_data_a = 16'b1111110010101000;
            14'h2669: o_data_a = 16'b1111110000010000;
            14'h266a: o_data_a = 16'b0000000000000100;
            14'h266b: o_data_a = 16'b1110001100001000;
            14'h266c: o_data_a = 16'b0000000000000101;
            14'h266d: o_data_a = 16'b1111110000010000;
            14'h266e: o_data_a = 16'b0000000000000000;
            14'h266f: o_data_a = 16'b1111110111101000;
            14'h2670: o_data_a = 16'b1110110010100000;
            14'h2671: o_data_a = 16'b1110001100001000;
            14'h2672: o_data_a = 16'b0000000000000000;
            14'h2673: o_data_a = 16'b1111110010101000;
            14'h2674: o_data_a = 16'b1111110000010000;
            14'h2675: o_data_a = 16'b0000000000000100;
            14'h2676: o_data_a = 16'b1111110000100000;
            14'h2677: o_data_a = 16'b1110001100001000;
            14'h2678: o_data_a = 16'b0000000000000000;
            14'h2679: o_data_a = 16'b1111110111001000;
            14'h267a: o_data_a = 16'b1111110010100000;
            14'h267b: o_data_a = 16'b1110101010001000;
            14'h267c: o_data_a = 16'b0000000000110110;
            14'h267d: o_data_a = 16'b1110101010000111;
            14'h267e: o_data_a = 16'b0100000000000000;
            14'h267f: o_data_a = 16'b1110110000010000;
            14'h2680: o_data_a = 16'b0000000000000000;
            14'h2681: o_data_a = 16'b1111110111101000;
            14'h2682: o_data_a = 16'b1110110010100000;
            14'h2683: o_data_a = 16'b1110001100001000;
            14'h2684: o_data_a = 16'b0000000000000000;
            14'h2685: o_data_a = 16'b1111110010101000;
            14'h2686: o_data_a = 16'b1111110000010000;
            14'h2687: o_data_a = 16'b0000000000010100;
            14'h2688: o_data_a = 16'b1110001100001000;
            14'h2689: o_data_a = 16'b0000000000000000;
            14'h268a: o_data_a = 16'b1111110111001000;
            14'h268b: o_data_a = 16'b1111110010100000;
            14'h268c: o_data_a = 16'b1110101010001000;
            14'h268d: o_data_a = 16'b0000000000000000;
            14'h268e: o_data_a = 16'b1111110010100000;
            14'h268f: o_data_a = 16'b1111110001001000;
            14'h2690: o_data_a = 16'b0000000000000000;
            14'h2691: o_data_a = 16'b1111110010101000;
            14'h2692: o_data_a = 16'b1111110000010000;
            14'h2693: o_data_a = 16'b0000000000010101;
            14'h2694: o_data_a = 16'b1110001100001000;
            14'h2695: o_data_a = 16'b0000000000100000;
            14'h2696: o_data_a = 16'b1110110000010000;
            14'h2697: o_data_a = 16'b0000000000000000;
            14'h2698: o_data_a = 16'b1111110111101000;
            14'h2699: o_data_a = 16'b1110110010100000;
            14'h269a: o_data_a = 16'b1110001100001000;
            14'h269b: o_data_a = 16'b0000000000000000;
            14'h269c: o_data_a = 16'b1111110010101000;
            14'h269d: o_data_a = 16'b1111110000010000;
            14'h269e: o_data_a = 16'b0000000000010110;
            14'h269f: o_data_a = 16'b1110001100001000;
            14'h26a0: o_data_a = 16'b0000000000000000;
            14'h26a1: o_data_a = 16'b1111110111001000;
            14'h26a2: o_data_a = 16'b1111110010100000;
            14'h26a3: o_data_a = 16'b1110101010001000;
            14'h26a4: o_data_a = 16'b0000000000000000;
            14'h26a5: o_data_a = 16'b1111110010101000;
            14'h26a6: o_data_a = 16'b1111110000010000;
            14'h26a7: o_data_a = 16'b0000000000010111;
            14'h26a8: o_data_a = 16'b1110001100001000;
            14'h26a9: o_data_a = 16'b0000000000000110;
            14'h26aa: o_data_a = 16'b1110110000010000;
            14'h26ab: o_data_a = 16'b0000000000000000;
            14'h26ac: o_data_a = 16'b1111110111101000;
            14'h26ad: o_data_a = 16'b1110110010100000;
            14'h26ae: o_data_a = 16'b1110001100001000;
            14'h26af: o_data_a = 16'b0000000000000001;
            14'h26b0: o_data_a = 16'b1110110000010000;
            14'h26b1: o_data_a = 16'b0000000000001101;
            14'h26b2: o_data_a = 16'b1110001100001000;
            14'h26b3: o_data_a = 16'b0110001000010001;
            14'h26b4: o_data_a = 16'b1110110000010000;
            14'h26b5: o_data_a = 16'b0000000000001110;
            14'h26b6: o_data_a = 16'b1110001100001000;
            14'h26b7: o_data_a = 16'b0010011010111011;
            14'h26b8: o_data_a = 16'b1110110000010000;
            14'h26b9: o_data_a = 16'b0000000001011111;
            14'h26ba: o_data_a = 16'b1110101010000111;
            14'h26bb: o_data_a = 16'b0000000000000000;
            14'h26bc: o_data_a = 16'b1111110010101000;
            14'h26bd: o_data_a = 16'b1111110000010000;
            14'h26be: o_data_a = 16'b0000000000011000;
            14'h26bf: o_data_a = 16'b1110001100001000;
            14'h26c0: o_data_a = 16'b0000000000000000;
            14'h26c1: o_data_a = 16'b1110110000010000;
            14'h26c2: o_data_a = 16'b0000000000001101;
            14'h26c3: o_data_a = 16'b1110001100001000;
            14'h26c4: o_data_a = 16'b0010011011101000;
            14'h26c5: o_data_a = 16'b1110110000010000;
            14'h26c6: o_data_a = 16'b0000000000001110;
            14'h26c7: o_data_a = 16'b1110001100001000;
            14'h26c8: o_data_a = 16'b0010011011001100;
            14'h26c9: o_data_a = 16'b1110110000010000;
            14'h26ca: o_data_a = 16'b0000000001011111;
            14'h26cb: o_data_a = 16'b1110101010000111;
            14'h26cc: o_data_a = 16'b0000000000000000;
            14'h26cd: o_data_a = 16'b1111110010101000;
            14'h26ce: o_data_a = 16'b1111110000010000;
            14'h26cf: o_data_a = 16'b0000000000000101;
            14'h26d0: o_data_a = 16'b1110001100001000;
            14'h26d1: o_data_a = 16'b0000000000000000;
            14'h26d2: o_data_a = 16'b1110110000010000;
            14'h26d3: o_data_a = 16'b0000000000001101;
            14'h26d4: o_data_a = 16'b1110001100001000;
            14'h26d5: o_data_a = 16'b0100100000011000;
            14'h26d6: o_data_a = 16'b1110110000010000;
            14'h26d7: o_data_a = 16'b0000000000001110;
            14'h26d8: o_data_a = 16'b1110001100001000;
            14'h26d9: o_data_a = 16'b0010011011011101;
            14'h26da: o_data_a = 16'b1110110000010000;
            14'h26db: o_data_a = 16'b0000000001011111;
            14'h26dc: o_data_a = 16'b1110101010000111;
            14'h26dd: o_data_a = 16'b0000000000000000;
            14'h26de: o_data_a = 16'b1111110010101000;
            14'h26df: o_data_a = 16'b1111110000010000;
            14'h26e0: o_data_a = 16'b0000000000000101;
            14'h26e1: o_data_a = 16'b1110001100001000;
            14'h26e2: o_data_a = 16'b0000000000000000;
            14'h26e3: o_data_a = 16'b1111110111001000;
            14'h26e4: o_data_a = 16'b1111110010100000;
            14'h26e5: o_data_a = 16'b1110101010001000;
            14'h26e6: o_data_a = 16'b0000000000110110;
            14'h26e7: o_data_a = 16'b1110101010000111;
            14'h26e8: o_data_a = 16'b0000000001111111;
            14'h26e9: o_data_a = 16'b1110110000010000;
            14'h26ea: o_data_a = 16'b0000000000000000;
            14'h26eb: o_data_a = 16'b1111110111101000;
            14'h26ec: o_data_a = 16'b1110110010100000;
            14'h26ed: o_data_a = 16'b1110001100001000;
            14'h26ee: o_data_a = 16'b0000000000000001;
            14'h26ef: o_data_a = 16'b1110110000010000;
            14'h26f0: o_data_a = 16'b0000000000001101;
            14'h26f1: o_data_a = 16'b1110001100001000;
            14'h26f2: o_data_a = 16'b0001011010110000;
            14'h26f3: o_data_a = 16'b1110110000010000;
            14'h26f4: o_data_a = 16'b0000000000001110;
            14'h26f5: o_data_a = 16'b1110001100001000;
            14'h26f6: o_data_a = 16'b0010011011111010;
            14'h26f7: o_data_a = 16'b1110110000010000;
            14'h26f8: o_data_a = 16'b0000000001011111;
            14'h26f9: o_data_a = 16'b1110101010000111;
            14'h26fa: o_data_a = 16'b0000000000000000;
            14'h26fb: o_data_a = 16'b1111110010101000;
            14'h26fc: o_data_a = 16'b1111110000010000;
            14'h26fd: o_data_a = 16'b0000000000011001;
            14'h26fe: o_data_a = 16'b1110001100001000;
            14'h26ff: o_data_a = 16'b0000000000000000;
            14'h2700: o_data_a = 16'b1111110111001000;
            14'h2701: o_data_a = 16'b1111110010100000;
            14'h2702: o_data_a = 16'b1110101010001000;
            14'h2703: o_data_a = 16'b0000000000111111;
            14'h2704: o_data_a = 16'b1110110000010000;
            14'h2705: o_data_a = 16'b0000000000000000;
            14'h2706: o_data_a = 16'b1111110111101000;
            14'h2707: o_data_a = 16'b1110110010100000;
            14'h2708: o_data_a = 16'b1110001100001000;
            14'h2709: o_data_a = 16'b0000000000111111;
            14'h270a: o_data_a = 16'b1110110000010000;
            14'h270b: o_data_a = 16'b0000000000000000;
            14'h270c: o_data_a = 16'b1111110111101000;
            14'h270d: o_data_a = 16'b1110110010100000;
            14'h270e: o_data_a = 16'b1110001100001000;
            14'h270f: o_data_a = 16'b0000000000111111;
            14'h2710: o_data_a = 16'b1110110000010000;
            14'h2711: o_data_a = 16'b0000000000000000;
            14'h2712: o_data_a = 16'b1111110111101000;
            14'h2713: o_data_a = 16'b1110110010100000;
            14'h2714: o_data_a = 16'b1110001100001000;
            14'h2715: o_data_a = 16'b0000000000111111;
            14'h2716: o_data_a = 16'b1110110000010000;
            14'h2717: o_data_a = 16'b0000000000000000;
            14'h2718: o_data_a = 16'b1111110111101000;
            14'h2719: o_data_a = 16'b1110110010100000;
            14'h271a: o_data_a = 16'b1110001100001000;
            14'h271b: o_data_a = 16'b0000000000111111;
            14'h271c: o_data_a = 16'b1110110000010000;
            14'h271d: o_data_a = 16'b0000000000000000;
            14'h271e: o_data_a = 16'b1111110111101000;
            14'h271f: o_data_a = 16'b1110110010100000;
            14'h2720: o_data_a = 16'b1110001100001000;
            14'h2721: o_data_a = 16'b0000000000111111;
            14'h2722: o_data_a = 16'b1110110000010000;
            14'h2723: o_data_a = 16'b0000000000000000;
            14'h2724: o_data_a = 16'b1111110111101000;
            14'h2725: o_data_a = 16'b1110110010100000;
            14'h2726: o_data_a = 16'b1110001100001000;
            14'h2727: o_data_a = 16'b0000000000111111;
            14'h2728: o_data_a = 16'b1110110000010000;
            14'h2729: o_data_a = 16'b0000000000000000;
            14'h272a: o_data_a = 16'b1111110111101000;
            14'h272b: o_data_a = 16'b1110110010100000;
            14'h272c: o_data_a = 16'b1110001100001000;
            14'h272d: o_data_a = 16'b0000000000111111;
            14'h272e: o_data_a = 16'b1110110000010000;
            14'h272f: o_data_a = 16'b0000000000000000;
            14'h2730: o_data_a = 16'b1111110111101000;
            14'h2731: o_data_a = 16'b1110110010100000;
            14'h2732: o_data_a = 16'b1110001100001000;
            14'h2733: o_data_a = 16'b0000000000111111;
            14'h2734: o_data_a = 16'b1110110000010000;
            14'h2735: o_data_a = 16'b0000000000000000;
            14'h2736: o_data_a = 16'b1111110111101000;
            14'h2737: o_data_a = 16'b1110110010100000;
            14'h2738: o_data_a = 16'b1110001100001000;
            14'h2739: o_data_a = 16'b0000000000000000;
            14'h273a: o_data_a = 16'b1111110111001000;
            14'h273b: o_data_a = 16'b1111110010100000;
            14'h273c: o_data_a = 16'b1110101010001000;
            14'h273d: o_data_a = 16'b0000000000000000;
            14'h273e: o_data_a = 16'b1111110111001000;
            14'h273f: o_data_a = 16'b1111110010100000;
            14'h2740: o_data_a = 16'b1110101010001000;
            14'h2741: o_data_a = 16'b0000000000001100;
            14'h2742: o_data_a = 16'b1110110000010000;
            14'h2743: o_data_a = 16'b0000000000001101;
            14'h2744: o_data_a = 16'b1110001100001000;
            14'h2745: o_data_a = 16'b0100010110110011;
            14'h2746: o_data_a = 16'b1110110000010000;
            14'h2747: o_data_a = 16'b0000000000001110;
            14'h2748: o_data_a = 16'b1110001100001000;
            14'h2749: o_data_a = 16'b0010011101001101;
            14'h274a: o_data_a = 16'b1110110000010000;
            14'h274b: o_data_a = 16'b0000000001011111;
            14'h274c: o_data_a = 16'b1110101010000111;
            14'h274d: o_data_a = 16'b0000000000000000;
            14'h274e: o_data_a = 16'b1111110010101000;
            14'h274f: o_data_a = 16'b1111110000010000;
            14'h2750: o_data_a = 16'b0000000000000101;
            14'h2751: o_data_a = 16'b1110001100001000;
            14'h2752: o_data_a = 16'b0000000000100000;
            14'h2753: o_data_a = 16'b1110110000010000;
            14'h2754: o_data_a = 16'b0000000000000000;
            14'h2755: o_data_a = 16'b1111110111101000;
            14'h2756: o_data_a = 16'b1110110010100000;
            14'h2757: o_data_a = 16'b1110001100001000;
            14'h2758: o_data_a = 16'b0000000000000000;
            14'h2759: o_data_a = 16'b1111110111001000;
            14'h275a: o_data_a = 16'b1111110010100000;
            14'h275b: o_data_a = 16'b1110101010001000;
            14'h275c: o_data_a = 16'b0000000000000000;
            14'h275d: o_data_a = 16'b1111110111001000;
            14'h275e: o_data_a = 16'b1111110010100000;
            14'h275f: o_data_a = 16'b1110101010001000;
            14'h2760: o_data_a = 16'b0000000000000000;
            14'h2761: o_data_a = 16'b1111110111001000;
            14'h2762: o_data_a = 16'b1111110010100000;
            14'h2763: o_data_a = 16'b1110101010001000;
            14'h2764: o_data_a = 16'b0000000000000000;
            14'h2765: o_data_a = 16'b1111110111001000;
            14'h2766: o_data_a = 16'b1111110010100000;
            14'h2767: o_data_a = 16'b1110101010001000;
            14'h2768: o_data_a = 16'b0000000000000000;
            14'h2769: o_data_a = 16'b1111110111001000;
            14'h276a: o_data_a = 16'b1111110010100000;
            14'h276b: o_data_a = 16'b1110101010001000;
            14'h276c: o_data_a = 16'b0000000000000000;
            14'h276d: o_data_a = 16'b1111110111001000;
            14'h276e: o_data_a = 16'b1111110010100000;
            14'h276f: o_data_a = 16'b1110101010001000;
            14'h2770: o_data_a = 16'b0000000000000000;
            14'h2771: o_data_a = 16'b1111110111001000;
            14'h2772: o_data_a = 16'b1111110010100000;
            14'h2773: o_data_a = 16'b1110101010001000;
            14'h2774: o_data_a = 16'b0000000000000000;
            14'h2775: o_data_a = 16'b1111110111001000;
            14'h2776: o_data_a = 16'b1111110010100000;
            14'h2777: o_data_a = 16'b1110101010001000;
            14'h2778: o_data_a = 16'b0000000000000000;
            14'h2779: o_data_a = 16'b1111110111001000;
            14'h277a: o_data_a = 16'b1111110010100000;
            14'h277b: o_data_a = 16'b1110101010001000;
            14'h277c: o_data_a = 16'b0000000000000000;
            14'h277d: o_data_a = 16'b1111110111001000;
            14'h277e: o_data_a = 16'b1111110010100000;
            14'h277f: o_data_a = 16'b1110101010001000;
            14'h2780: o_data_a = 16'b0000000000000000;
            14'h2781: o_data_a = 16'b1111110111001000;
            14'h2782: o_data_a = 16'b1111110010100000;
            14'h2783: o_data_a = 16'b1110101010001000;
            14'h2784: o_data_a = 16'b0000000000001100;
            14'h2785: o_data_a = 16'b1110110000010000;
            14'h2786: o_data_a = 16'b0000000000001101;
            14'h2787: o_data_a = 16'b1110001100001000;
            14'h2788: o_data_a = 16'b0100010110110011;
            14'h2789: o_data_a = 16'b1110110000010000;
            14'h278a: o_data_a = 16'b0000000000001110;
            14'h278b: o_data_a = 16'b1110001100001000;
            14'h278c: o_data_a = 16'b0010011110010000;
            14'h278d: o_data_a = 16'b1110110000010000;
            14'h278e: o_data_a = 16'b0000000001011111;
            14'h278f: o_data_a = 16'b1110101010000111;
            14'h2790: o_data_a = 16'b0000000000000000;
            14'h2791: o_data_a = 16'b1111110010101000;
            14'h2792: o_data_a = 16'b1111110000010000;
            14'h2793: o_data_a = 16'b0000000000000101;
            14'h2794: o_data_a = 16'b1110001100001000;
            14'h2795: o_data_a = 16'b0000000000100001;
            14'h2796: o_data_a = 16'b1110110000010000;
            14'h2797: o_data_a = 16'b0000000000000000;
            14'h2798: o_data_a = 16'b1111110111101000;
            14'h2799: o_data_a = 16'b1110110010100000;
            14'h279a: o_data_a = 16'b1110001100001000;
            14'h279b: o_data_a = 16'b0000000000001100;
            14'h279c: o_data_a = 16'b1110110000010000;
            14'h279d: o_data_a = 16'b0000000000000000;
            14'h279e: o_data_a = 16'b1111110111101000;
            14'h279f: o_data_a = 16'b1110110010100000;
            14'h27a0: o_data_a = 16'b1110001100001000;
            14'h27a1: o_data_a = 16'b0000000000011110;
            14'h27a2: o_data_a = 16'b1110110000010000;
            14'h27a3: o_data_a = 16'b0000000000000000;
            14'h27a4: o_data_a = 16'b1111110111101000;
            14'h27a5: o_data_a = 16'b1110110010100000;
            14'h27a6: o_data_a = 16'b1110001100001000;
            14'h27a7: o_data_a = 16'b0000000000011110;
            14'h27a8: o_data_a = 16'b1110110000010000;
            14'h27a9: o_data_a = 16'b0000000000000000;
            14'h27aa: o_data_a = 16'b1111110111101000;
            14'h27ab: o_data_a = 16'b1110110010100000;
            14'h27ac: o_data_a = 16'b1110001100001000;
            14'h27ad: o_data_a = 16'b0000000000011110;
            14'h27ae: o_data_a = 16'b1110110000010000;
            14'h27af: o_data_a = 16'b0000000000000000;
            14'h27b0: o_data_a = 16'b1111110111101000;
            14'h27b1: o_data_a = 16'b1110110010100000;
            14'h27b2: o_data_a = 16'b1110001100001000;
            14'h27b3: o_data_a = 16'b0000000000001100;
            14'h27b4: o_data_a = 16'b1110110000010000;
            14'h27b5: o_data_a = 16'b0000000000000000;
            14'h27b6: o_data_a = 16'b1111110111101000;
            14'h27b7: o_data_a = 16'b1110110010100000;
            14'h27b8: o_data_a = 16'b1110001100001000;
            14'h27b9: o_data_a = 16'b0000000000001100;
            14'h27ba: o_data_a = 16'b1110110000010000;
            14'h27bb: o_data_a = 16'b0000000000000000;
            14'h27bc: o_data_a = 16'b1111110111101000;
            14'h27bd: o_data_a = 16'b1110110010100000;
            14'h27be: o_data_a = 16'b1110001100001000;
            14'h27bf: o_data_a = 16'b0000000000000000;
            14'h27c0: o_data_a = 16'b1111110111001000;
            14'h27c1: o_data_a = 16'b1111110010100000;
            14'h27c2: o_data_a = 16'b1110101010001000;
            14'h27c3: o_data_a = 16'b0000000000001100;
            14'h27c4: o_data_a = 16'b1110110000010000;
            14'h27c5: o_data_a = 16'b0000000000000000;
            14'h27c6: o_data_a = 16'b1111110111101000;
            14'h27c7: o_data_a = 16'b1110110010100000;
            14'h27c8: o_data_a = 16'b1110001100001000;
            14'h27c9: o_data_a = 16'b0000000000001100;
            14'h27ca: o_data_a = 16'b1110110000010000;
            14'h27cb: o_data_a = 16'b0000000000000000;
            14'h27cc: o_data_a = 16'b1111110111101000;
            14'h27cd: o_data_a = 16'b1110110010100000;
            14'h27ce: o_data_a = 16'b1110001100001000;
            14'h27cf: o_data_a = 16'b0000000000000000;
            14'h27d0: o_data_a = 16'b1111110111001000;
            14'h27d1: o_data_a = 16'b1111110010100000;
            14'h27d2: o_data_a = 16'b1110101010001000;
            14'h27d3: o_data_a = 16'b0000000000000000;
            14'h27d4: o_data_a = 16'b1111110111001000;
            14'h27d5: o_data_a = 16'b1111110010100000;
            14'h27d6: o_data_a = 16'b1110101010001000;
            14'h27d7: o_data_a = 16'b0000000000001100;
            14'h27d8: o_data_a = 16'b1110110000010000;
            14'h27d9: o_data_a = 16'b0000000000001101;
            14'h27da: o_data_a = 16'b1110001100001000;
            14'h27db: o_data_a = 16'b0100010110110011;
            14'h27dc: o_data_a = 16'b1110110000010000;
            14'h27dd: o_data_a = 16'b0000000000001110;
            14'h27de: o_data_a = 16'b1110001100001000;
            14'h27df: o_data_a = 16'b0010011111100011;
            14'h27e0: o_data_a = 16'b1110110000010000;
            14'h27e1: o_data_a = 16'b0000000001011111;
            14'h27e2: o_data_a = 16'b1110101010000111;
            14'h27e3: o_data_a = 16'b0000000000000000;
            14'h27e4: o_data_a = 16'b1111110010101000;
            14'h27e5: o_data_a = 16'b1111110000010000;
            14'h27e6: o_data_a = 16'b0000000000000101;
            14'h27e7: o_data_a = 16'b1110001100001000;
            14'h27e8: o_data_a = 16'b0000000000100010;
            14'h27e9: o_data_a = 16'b1110110000010000;
            14'h27ea: o_data_a = 16'b0000000000000000;
            14'h27eb: o_data_a = 16'b1111110111101000;
            14'h27ec: o_data_a = 16'b1110110010100000;
            14'h27ed: o_data_a = 16'b1110001100001000;
            14'h27ee: o_data_a = 16'b0000000000110110;
            14'h27ef: o_data_a = 16'b1110110000010000;
            14'h27f0: o_data_a = 16'b0000000000000000;
            14'h27f1: o_data_a = 16'b1111110111101000;
            14'h27f2: o_data_a = 16'b1110110010100000;
            14'h27f3: o_data_a = 16'b1110001100001000;
            14'h27f4: o_data_a = 16'b0000000000110110;
            14'h27f5: o_data_a = 16'b1110110000010000;
            14'h27f6: o_data_a = 16'b0000000000000000;
            14'h27f7: o_data_a = 16'b1111110111101000;
            14'h27f8: o_data_a = 16'b1110110010100000;
            14'h27f9: o_data_a = 16'b1110001100001000;
            14'h27fa: o_data_a = 16'b0000000000010100;
            14'h27fb: o_data_a = 16'b1110110000010000;
            14'h27fc: o_data_a = 16'b0000000000000000;
            14'h27fd: o_data_a = 16'b1111110111101000;
            14'h27fe: o_data_a = 16'b1110110010100000;
            14'h27ff: o_data_a = 16'b1110001100001000;
            14'h2800: o_data_a = 16'b0000000000000000;
            14'h2801: o_data_a = 16'b1111110111001000;
            14'h2802: o_data_a = 16'b1111110010100000;
            14'h2803: o_data_a = 16'b1110101010001000;
            14'h2804: o_data_a = 16'b0000000000000000;
            14'h2805: o_data_a = 16'b1111110111001000;
            14'h2806: o_data_a = 16'b1111110010100000;
            14'h2807: o_data_a = 16'b1110101010001000;
            14'h2808: o_data_a = 16'b0000000000000000;
            14'h2809: o_data_a = 16'b1111110111001000;
            14'h280a: o_data_a = 16'b1111110010100000;
            14'h280b: o_data_a = 16'b1110101010001000;
            14'h280c: o_data_a = 16'b0000000000000000;
            14'h280d: o_data_a = 16'b1111110111001000;
            14'h280e: o_data_a = 16'b1111110010100000;
            14'h280f: o_data_a = 16'b1110101010001000;
            14'h2810: o_data_a = 16'b0000000000000000;
            14'h2811: o_data_a = 16'b1111110111001000;
            14'h2812: o_data_a = 16'b1111110010100000;
            14'h2813: o_data_a = 16'b1110101010001000;
            14'h2814: o_data_a = 16'b0000000000000000;
            14'h2815: o_data_a = 16'b1111110111001000;
            14'h2816: o_data_a = 16'b1111110010100000;
            14'h2817: o_data_a = 16'b1110101010001000;
            14'h2818: o_data_a = 16'b0000000000000000;
            14'h2819: o_data_a = 16'b1111110111001000;
            14'h281a: o_data_a = 16'b1111110010100000;
            14'h281b: o_data_a = 16'b1110101010001000;
            14'h281c: o_data_a = 16'b0000000000000000;
            14'h281d: o_data_a = 16'b1111110111001000;
            14'h281e: o_data_a = 16'b1111110010100000;
            14'h281f: o_data_a = 16'b1110101010001000;
            14'h2820: o_data_a = 16'b0000000000001100;
            14'h2821: o_data_a = 16'b1110110000010000;
            14'h2822: o_data_a = 16'b0000000000001101;
            14'h2823: o_data_a = 16'b1110001100001000;
            14'h2824: o_data_a = 16'b0100010110110011;
            14'h2825: o_data_a = 16'b1110110000010000;
            14'h2826: o_data_a = 16'b0000000000001110;
            14'h2827: o_data_a = 16'b1110001100001000;
            14'h2828: o_data_a = 16'b0010100000101100;
            14'h2829: o_data_a = 16'b1110110000010000;
            14'h282a: o_data_a = 16'b0000000001011111;
            14'h282b: o_data_a = 16'b1110101010000111;
            14'h282c: o_data_a = 16'b0000000000000000;
            14'h282d: o_data_a = 16'b1111110010101000;
            14'h282e: o_data_a = 16'b1111110000010000;
            14'h282f: o_data_a = 16'b0000000000000101;
            14'h2830: o_data_a = 16'b1110001100001000;
            14'h2831: o_data_a = 16'b0000000000100011;
            14'h2832: o_data_a = 16'b1110110000010000;
            14'h2833: o_data_a = 16'b0000000000000000;
            14'h2834: o_data_a = 16'b1111110111101000;
            14'h2835: o_data_a = 16'b1110110010100000;
            14'h2836: o_data_a = 16'b1110001100001000;
            14'h2837: o_data_a = 16'b0000000000000000;
            14'h2838: o_data_a = 16'b1111110111001000;
            14'h2839: o_data_a = 16'b1111110010100000;
            14'h283a: o_data_a = 16'b1110101010001000;
            14'h283b: o_data_a = 16'b0000000000010010;
            14'h283c: o_data_a = 16'b1110110000010000;
            14'h283d: o_data_a = 16'b0000000000000000;
            14'h283e: o_data_a = 16'b1111110111101000;
            14'h283f: o_data_a = 16'b1110110010100000;
            14'h2840: o_data_a = 16'b1110001100001000;
            14'h2841: o_data_a = 16'b0000000000010010;
            14'h2842: o_data_a = 16'b1110110000010000;
            14'h2843: o_data_a = 16'b0000000000000000;
            14'h2844: o_data_a = 16'b1111110111101000;
            14'h2845: o_data_a = 16'b1110110010100000;
            14'h2846: o_data_a = 16'b1110001100001000;
            14'h2847: o_data_a = 16'b0000000000111111;
            14'h2848: o_data_a = 16'b1110110000010000;
            14'h2849: o_data_a = 16'b0000000000000000;
            14'h284a: o_data_a = 16'b1111110111101000;
            14'h284b: o_data_a = 16'b1110110010100000;
            14'h284c: o_data_a = 16'b1110001100001000;
            14'h284d: o_data_a = 16'b0000000000010010;
            14'h284e: o_data_a = 16'b1110110000010000;
            14'h284f: o_data_a = 16'b0000000000000000;
            14'h2850: o_data_a = 16'b1111110111101000;
            14'h2851: o_data_a = 16'b1110110010100000;
            14'h2852: o_data_a = 16'b1110001100001000;
            14'h2853: o_data_a = 16'b0000000000010010;
            14'h2854: o_data_a = 16'b1110110000010000;
            14'h2855: o_data_a = 16'b0000000000000000;
            14'h2856: o_data_a = 16'b1111110111101000;
            14'h2857: o_data_a = 16'b1110110010100000;
            14'h2858: o_data_a = 16'b1110001100001000;
            14'h2859: o_data_a = 16'b0000000000111111;
            14'h285a: o_data_a = 16'b1110110000010000;
            14'h285b: o_data_a = 16'b0000000000000000;
            14'h285c: o_data_a = 16'b1111110111101000;
            14'h285d: o_data_a = 16'b1110110010100000;
            14'h285e: o_data_a = 16'b1110001100001000;
            14'h285f: o_data_a = 16'b0000000000010010;
            14'h2860: o_data_a = 16'b1110110000010000;
            14'h2861: o_data_a = 16'b0000000000000000;
            14'h2862: o_data_a = 16'b1111110111101000;
            14'h2863: o_data_a = 16'b1110110010100000;
            14'h2864: o_data_a = 16'b1110001100001000;
            14'h2865: o_data_a = 16'b0000000000010010;
            14'h2866: o_data_a = 16'b1110110000010000;
            14'h2867: o_data_a = 16'b0000000000000000;
            14'h2868: o_data_a = 16'b1111110111101000;
            14'h2869: o_data_a = 16'b1110110010100000;
            14'h286a: o_data_a = 16'b1110001100001000;
            14'h286b: o_data_a = 16'b0000000000000000;
            14'h286c: o_data_a = 16'b1111110111001000;
            14'h286d: o_data_a = 16'b1111110010100000;
            14'h286e: o_data_a = 16'b1110101010001000;
            14'h286f: o_data_a = 16'b0000000000000000;
            14'h2870: o_data_a = 16'b1111110111001000;
            14'h2871: o_data_a = 16'b1111110010100000;
            14'h2872: o_data_a = 16'b1110101010001000;
            14'h2873: o_data_a = 16'b0000000000001100;
            14'h2874: o_data_a = 16'b1110110000010000;
            14'h2875: o_data_a = 16'b0000000000001101;
            14'h2876: o_data_a = 16'b1110001100001000;
            14'h2877: o_data_a = 16'b0100010110110011;
            14'h2878: o_data_a = 16'b1110110000010000;
            14'h2879: o_data_a = 16'b0000000000001110;
            14'h287a: o_data_a = 16'b1110001100001000;
            14'h287b: o_data_a = 16'b0010100001111111;
            14'h287c: o_data_a = 16'b1110110000010000;
            14'h287d: o_data_a = 16'b0000000001011111;
            14'h287e: o_data_a = 16'b1110101010000111;
            14'h287f: o_data_a = 16'b0000000000000000;
            14'h2880: o_data_a = 16'b1111110010101000;
            14'h2881: o_data_a = 16'b1111110000010000;
            14'h2882: o_data_a = 16'b0000000000000101;
            14'h2883: o_data_a = 16'b1110001100001000;
            14'h2884: o_data_a = 16'b0000000000100100;
            14'h2885: o_data_a = 16'b1110110000010000;
            14'h2886: o_data_a = 16'b0000000000000000;
            14'h2887: o_data_a = 16'b1111110111101000;
            14'h2888: o_data_a = 16'b1110110010100000;
            14'h2889: o_data_a = 16'b1110001100001000;
            14'h288a: o_data_a = 16'b0000000000001100;
            14'h288b: o_data_a = 16'b1110110000010000;
            14'h288c: o_data_a = 16'b0000000000000000;
            14'h288d: o_data_a = 16'b1111110111101000;
            14'h288e: o_data_a = 16'b1110110010100000;
            14'h288f: o_data_a = 16'b1110001100001000;
            14'h2890: o_data_a = 16'b0000000000011110;
            14'h2891: o_data_a = 16'b1110110000010000;
            14'h2892: o_data_a = 16'b0000000000000000;
            14'h2893: o_data_a = 16'b1111110111101000;
            14'h2894: o_data_a = 16'b1110110010100000;
            14'h2895: o_data_a = 16'b1110001100001000;
            14'h2896: o_data_a = 16'b0000000000110011;
            14'h2897: o_data_a = 16'b1110110000010000;
            14'h2898: o_data_a = 16'b0000000000000000;
            14'h2899: o_data_a = 16'b1111110111101000;
            14'h289a: o_data_a = 16'b1110110010100000;
            14'h289b: o_data_a = 16'b1110001100001000;
            14'h289c: o_data_a = 16'b0000000000000011;
            14'h289d: o_data_a = 16'b1110110000010000;
            14'h289e: o_data_a = 16'b0000000000000000;
            14'h289f: o_data_a = 16'b1111110111101000;
            14'h28a0: o_data_a = 16'b1110110010100000;
            14'h28a1: o_data_a = 16'b1110001100001000;
            14'h28a2: o_data_a = 16'b0000000000011110;
            14'h28a3: o_data_a = 16'b1110110000010000;
            14'h28a4: o_data_a = 16'b0000000000000000;
            14'h28a5: o_data_a = 16'b1111110111101000;
            14'h28a6: o_data_a = 16'b1110110010100000;
            14'h28a7: o_data_a = 16'b1110001100001000;
            14'h28a8: o_data_a = 16'b0000000000110000;
            14'h28a9: o_data_a = 16'b1110110000010000;
            14'h28aa: o_data_a = 16'b0000000000000000;
            14'h28ab: o_data_a = 16'b1111110111101000;
            14'h28ac: o_data_a = 16'b1110110010100000;
            14'h28ad: o_data_a = 16'b1110001100001000;
            14'h28ae: o_data_a = 16'b0000000000110011;
            14'h28af: o_data_a = 16'b1110110000010000;
            14'h28b0: o_data_a = 16'b0000000000000000;
            14'h28b1: o_data_a = 16'b1111110111101000;
            14'h28b2: o_data_a = 16'b1110110010100000;
            14'h28b3: o_data_a = 16'b1110001100001000;
            14'h28b4: o_data_a = 16'b0000000000011110;
            14'h28b5: o_data_a = 16'b1110110000010000;
            14'h28b6: o_data_a = 16'b0000000000000000;
            14'h28b7: o_data_a = 16'b1111110111101000;
            14'h28b8: o_data_a = 16'b1110110010100000;
            14'h28b9: o_data_a = 16'b1110001100001000;
            14'h28ba: o_data_a = 16'b0000000000001100;
            14'h28bb: o_data_a = 16'b1110110000010000;
            14'h28bc: o_data_a = 16'b0000000000000000;
            14'h28bd: o_data_a = 16'b1111110111101000;
            14'h28be: o_data_a = 16'b1110110010100000;
            14'h28bf: o_data_a = 16'b1110001100001000;
            14'h28c0: o_data_a = 16'b0000000000001100;
            14'h28c1: o_data_a = 16'b1110110000010000;
            14'h28c2: o_data_a = 16'b0000000000000000;
            14'h28c3: o_data_a = 16'b1111110111101000;
            14'h28c4: o_data_a = 16'b1110110010100000;
            14'h28c5: o_data_a = 16'b1110001100001000;
            14'h28c6: o_data_a = 16'b0000000000000000;
            14'h28c7: o_data_a = 16'b1111110111001000;
            14'h28c8: o_data_a = 16'b1111110010100000;
            14'h28c9: o_data_a = 16'b1110101010001000;
            14'h28ca: o_data_a = 16'b0000000000001100;
            14'h28cb: o_data_a = 16'b1110110000010000;
            14'h28cc: o_data_a = 16'b0000000000001101;
            14'h28cd: o_data_a = 16'b1110001100001000;
            14'h28ce: o_data_a = 16'b0100010110110011;
            14'h28cf: o_data_a = 16'b1110110000010000;
            14'h28d0: o_data_a = 16'b0000000000001110;
            14'h28d1: o_data_a = 16'b1110001100001000;
            14'h28d2: o_data_a = 16'b0010100011010110;
            14'h28d3: o_data_a = 16'b1110110000010000;
            14'h28d4: o_data_a = 16'b0000000001011111;
            14'h28d5: o_data_a = 16'b1110101010000111;
            14'h28d6: o_data_a = 16'b0000000000000000;
            14'h28d7: o_data_a = 16'b1111110010101000;
            14'h28d8: o_data_a = 16'b1111110000010000;
            14'h28d9: o_data_a = 16'b0000000000000101;
            14'h28da: o_data_a = 16'b1110001100001000;
            14'h28db: o_data_a = 16'b0000000000100101;
            14'h28dc: o_data_a = 16'b1110110000010000;
            14'h28dd: o_data_a = 16'b0000000000000000;
            14'h28de: o_data_a = 16'b1111110111101000;
            14'h28df: o_data_a = 16'b1110110010100000;
            14'h28e0: o_data_a = 16'b1110001100001000;
            14'h28e1: o_data_a = 16'b0000000000000000;
            14'h28e2: o_data_a = 16'b1111110111001000;
            14'h28e3: o_data_a = 16'b1111110010100000;
            14'h28e4: o_data_a = 16'b1110101010001000;
            14'h28e5: o_data_a = 16'b0000000000000000;
            14'h28e6: o_data_a = 16'b1111110111001000;
            14'h28e7: o_data_a = 16'b1111110010100000;
            14'h28e8: o_data_a = 16'b1110101010001000;
            14'h28e9: o_data_a = 16'b0000000000100011;
            14'h28ea: o_data_a = 16'b1110110000010000;
            14'h28eb: o_data_a = 16'b0000000000000000;
            14'h28ec: o_data_a = 16'b1111110111101000;
            14'h28ed: o_data_a = 16'b1110110010100000;
            14'h28ee: o_data_a = 16'b1110001100001000;
            14'h28ef: o_data_a = 16'b0000000000110011;
            14'h28f0: o_data_a = 16'b1110110000010000;
            14'h28f1: o_data_a = 16'b0000000000000000;
            14'h28f2: o_data_a = 16'b1111110111101000;
            14'h28f3: o_data_a = 16'b1110110010100000;
            14'h28f4: o_data_a = 16'b1110001100001000;
            14'h28f5: o_data_a = 16'b0000000000011000;
            14'h28f6: o_data_a = 16'b1110110000010000;
            14'h28f7: o_data_a = 16'b0000000000000000;
            14'h28f8: o_data_a = 16'b1111110111101000;
            14'h28f9: o_data_a = 16'b1110110010100000;
            14'h28fa: o_data_a = 16'b1110001100001000;
            14'h28fb: o_data_a = 16'b0000000000001100;
            14'h28fc: o_data_a = 16'b1110110000010000;
            14'h28fd: o_data_a = 16'b0000000000000000;
            14'h28fe: o_data_a = 16'b1111110111101000;
            14'h28ff: o_data_a = 16'b1110110010100000;
            14'h2900: o_data_a = 16'b1110001100001000;
            14'h2901: o_data_a = 16'b0000000000000110;
            14'h2902: o_data_a = 16'b1110110000010000;
            14'h2903: o_data_a = 16'b0000000000000000;
            14'h2904: o_data_a = 16'b1111110111101000;
            14'h2905: o_data_a = 16'b1110110010100000;
            14'h2906: o_data_a = 16'b1110001100001000;
            14'h2907: o_data_a = 16'b0000000000110011;
            14'h2908: o_data_a = 16'b1110110000010000;
            14'h2909: o_data_a = 16'b0000000000000000;
            14'h290a: o_data_a = 16'b1111110111101000;
            14'h290b: o_data_a = 16'b1110110010100000;
            14'h290c: o_data_a = 16'b1110001100001000;
            14'h290d: o_data_a = 16'b0000000000110001;
            14'h290e: o_data_a = 16'b1110110000010000;
            14'h290f: o_data_a = 16'b0000000000000000;
            14'h2910: o_data_a = 16'b1111110111101000;
            14'h2911: o_data_a = 16'b1110110010100000;
            14'h2912: o_data_a = 16'b1110001100001000;
            14'h2913: o_data_a = 16'b0000000000000000;
            14'h2914: o_data_a = 16'b1111110111001000;
            14'h2915: o_data_a = 16'b1111110010100000;
            14'h2916: o_data_a = 16'b1110101010001000;
            14'h2917: o_data_a = 16'b0000000000000000;
            14'h2918: o_data_a = 16'b1111110111001000;
            14'h2919: o_data_a = 16'b1111110010100000;
            14'h291a: o_data_a = 16'b1110101010001000;
            14'h291b: o_data_a = 16'b0000000000001100;
            14'h291c: o_data_a = 16'b1110110000010000;
            14'h291d: o_data_a = 16'b0000000000001101;
            14'h291e: o_data_a = 16'b1110001100001000;
            14'h291f: o_data_a = 16'b0100010110110011;
            14'h2920: o_data_a = 16'b1110110000010000;
            14'h2921: o_data_a = 16'b0000000000001110;
            14'h2922: o_data_a = 16'b1110001100001000;
            14'h2923: o_data_a = 16'b0010100100100111;
            14'h2924: o_data_a = 16'b1110110000010000;
            14'h2925: o_data_a = 16'b0000000001011111;
            14'h2926: o_data_a = 16'b1110101010000111;
            14'h2927: o_data_a = 16'b0000000000000000;
            14'h2928: o_data_a = 16'b1111110010101000;
            14'h2929: o_data_a = 16'b1111110000010000;
            14'h292a: o_data_a = 16'b0000000000000101;
            14'h292b: o_data_a = 16'b1110001100001000;
            14'h292c: o_data_a = 16'b0000000000100110;
            14'h292d: o_data_a = 16'b1110110000010000;
            14'h292e: o_data_a = 16'b0000000000000000;
            14'h292f: o_data_a = 16'b1111110111101000;
            14'h2930: o_data_a = 16'b1110110010100000;
            14'h2931: o_data_a = 16'b1110001100001000;
            14'h2932: o_data_a = 16'b0000000000001100;
            14'h2933: o_data_a = 16'b1110110000010000;
            14'h2934: o_data_a = 16'b0000000000000000;
            14'h2935: o_data_a = 16'b1111110111101000;
            14'h2936: o_data_a = 16'b1110110010100000;
            14'h2937: o_data_a = 16'b1110001100001000;
            14'h2938: o_data_a = 16'b0000000000011110;
            14'h2939: o_data_a = 16'b1110110000010000;
            14'h293a: o_data_a = 16'b0000000000000000;
            14'h293b: o_data_a = 16'b1111110111101000;
            14'h293c: o_data_a = 16'b1110110010100000;
            14'h293d: o_data_a = 16'b1110001100001000;
            14'h293e: o_data_a = 16'b0000000000011110;
            14'h293f: o_data_a = 16'b1110110000010000;
            14'h2940: o_data_a = 16'b0000000000000000;
            14'h2941: o_data_a = 16'b1111110111101000;
            14'h2942: o_data_a = 16'b1110110010100000;
            14'h2943: o_data_a = 16'b1110001100001000;
            14'h2944: o_data_a = 16'b0000000000001100;
            14'h2945: o_data_a = 16'b1110110000010000;
            14'h2946: o_data_a = 16'b0000000000000000;
            14'h2947: o_data_a = 16'b1111110111101000;
            14'h2948: o_data_a = 16'b1110110010100000;
            14'h2949: o_data_a = 16'b1110001100001000;
            14'h294a: o_data_a = 16'b0000000000110110;
            14'h294b: o_data_a = 16'b1110110000010000;
            14'h294c: o_data_a = 16'b0000000000000000;
            14'h294d: o_data_a = 16'b1111110111101000;
            14'h294e: o_data_a = 16'b1110110010100000;
            14'h294f: o_data_a = 16'b1110001100001000;
            14'h2950: o_data_a = 16'b0000000000011011;
            14'h2951: o_data_a = 16'b1110110000010000;
            14'h2952: o_data_a = 16'b0000000000000000;
            14'h2953: o_data_a = 16'b1111110111101000;
            14'h2954: o_data_a = 16'b1110110010100000;
            14'h2955: o_data_a = 16'b1110001100001000;
            14'h2956: o_data_a = 16'b0000000000011011;
            14'h2957: o_data_a = 16'b1110110000010000;
            14'h2958: o_data_a = 16'b0000000000000000;
            14'h2959: o_data_a = 16'b1111110111101000;
            14'h295a: o_data_a = 16'b1110110010100000;
            14'h295b: o_data_a = 16'b1110001100001000;
            14'h295c: o_data_a = 16'b0000000000011011;
            14'h295d: o_data_a = 16'b1110110000010000;
            14'h295e: o_data_a = 16'b0000000000000000;
            14'h295f: o_data_a = 16'b1111110111101000;
            14'h2960: o_data_a = 16'b1110110010100000;
            14'h2961: o_data_a = 16'b1110001100001000;
            14'h2962: o_data_a = 16'b0000000000110110;
            14'h2963: o_data_a = 16'b1110110000010000;
            14'h2964: o_data_a = 16'b0000000000000000;
            14'h2965: o_data_a = 16'b1111110111101000;
            14'h2966: o_data_a = 16'b1110110010100000;
            14'h2967: o_data_a = 16'b1110001100001000;
            14'h2968: o_data_a = 16'b0000000000000000;
            14'h2969: o_data_a = 16'b1111110111001000;
            14'h296a: o_data_a = 16'b1111110010100000;
            14'h296b: o_data_a = 16'b1110101010001000;
            14'h296c: o_data_a = 16'b0000000000000000;
            14'h296d: o_data_a = 16'b1111110111001000;
            14'h296e: o_data_a = 16'b1111110010100000;
            14'h296f: o_data_a = 16'b1110101010001000;
            14'h2970: o_data_a = 16'b0000000000001100;
            14'h2971: o_data_a = 16'b1110110000010000;
            14'h2972: o_data_a = 16'b0000000000001101;
            14'h2973: o_data_a = 16'b1110001100001000;
            14'h2974: o_data_a = 16'b0100010110110011;
            14'h2975: o_data_a = 16'b1110110000010000;
            14'h2976: o_data_a = 16'b0000000000001110;
            14'h2977: o_data_a = 16'b1110001100001000;
            14'h2978: o_data_a = 16'b0010100101111100;
            14'h2979: o_data_a = 16'b1110110000010000;
            14'h297a: o_data_a = 16'b0000000001011111;
            14'h297b: o_data_a = 16'b1110101010000111;
            14'h297c: o_data_a = 16'b0000000000000000;
            14'h297d: o_data_a = 16'b1111110010101000;
            14'h297e: o_data_a = 16'b1111110000010000;
            14'h297f: o_data_a = 16'b0000000000000101;
            14'h2980: o_data_a = 16'b1110001100001000;
            14'h2981: o_data_a = 16'b0000000000100111;
            14'h2982: o_data_a = 16'b1110110000010000;
            14'h2983: o_data_a = 16'b0000000000000000;
            14'h2984: o_data_a = 16'b1111110111101000;
            14'h2985: o_data_a = 16'b1110110010100000;
            14'h2986: o_data_a = 16'b1110001100001000;
            14'h2987: o_data_a = 16'b0000000000001100;
            14'h2988: o_data_a = 16'b1110110000010000;
            14'h2989: o_data_a = 16'b0000000000000000;
            14'h298a: o_data_a = 16'b1111110111101000;
            14'h298b: o_data_a = 16'b1110110010100000;
            14'h298c: o_data_a = 16'b1110001100001000;
            14'h298d: o_data_a = 16'b0000000000001100;
            14'h298e: o_data_a = 16'b1110110000010000;
            14'h298f: o_data_a = 16'b0000000000000000;
            14'h2990: o_data_a = 16'b1111110111101000;
            14'h2991: o_data_a = 16'b1110110010100000;
            14'h2992: o_data_a = 16'b1110001100001000;
            14'h2993: o_data_a = 16'b0000000000000110;
            14'h2994: o_data_a = 16'b1110110000010000;
            14'h2995: o_data_a = 16'b0000000000000000;
            14'h2996: o_data_a = 16'b1111110111101000;
            14'h2997: o_data_a = 16'b1110110010100000;
            14'h2998: o_data_a = 16'b1110001100001000;
            14'h2999: o_data_a = 16'b0000000000000000;
            14'h299a: o_data_a = 16'b1111110111001000;
            14'h299b: o_data_a = 16'b1111110010100000;
            14'h299c: o_data_a = 16'b1110101010001000;
            14'h299d: o_data_a = 16'b0000000000000000;
            14'h299e: o_data_a = 16'b1111110111001000;
            14'h299f: o_data_a = 16'b1111110010100000;
            14'h29a0: o_data_a = 16'b1110101010001000;
            14'h29a1: o_data_a = 16'b0000000000000000;
            14'h29a2: o_data_a = 16'b1111110111001000;
            14'h29a3: o_data_a = 16'b1111110010100000;
            14'h29a4: o_data_a = 16'b1110101010001000;
            14'h29a5: o_data_a = 16'b0000000000000000;
            14'h29a6: o_data_a = 16'b1111110111001000;
            14'h29a7: o_data_a = 16'b1111110010100000;
            14'h29a8: o_data_a = 16'b1110101010001000;
            14'h29a9: o_data_a = 16'b0000000000000000;
            14'h29aa: o_data_a = 16'b1111110111001000;
            14'h29ab: o_data_a = 16'b1111110010100000;
            14'h29ac: o_data_a = 16'b1110101010001000;
            14'h29ad: o_data_a = 16'b0000000000000000;
            14'h29ae: o_data_a = 16'b1111110111001000;
            14'h29af: o_data_a = 16'b1111110010100000;
            14'h29b0: o_data_a = 16'b1110101010001000;
            14'h29b1: o_data_a = 16'b0000000000000000;
            14'h29b2: o_data_a = 16'b1111110111001000;
            14'h29b3: o_data_a = 16'b1111110010100000;
            14'h29b4: o_data_a = 16'b1110101010001000;
            14'h29b5: o_data_a = 16'b0000000000000000;
            14'h29b6: o_data_a = 16'b1111110111001000;
            14'h29b7: o_data_a = 16'b1111110010100000;
            14'h29b8: o_data_a = 16'b1110101010001000;
            14'h29b9: o_data_a = 16'b0000000000001100;
            14'h29ba: o_data_a = 16'b1110110000010000;
            14'h29bb: o_data_a = 16'b0000000000001101;
            14'h29bc: o_data_a = 16'b1110001100001000;
            14'h29bd: o_data_a = 16'b0100010110110011;
            14'h29be: o_data_a = 16'b1110110000010000;
            14'h29bf: o_data_a = 16'b0000000000001110;
            14'h29c0: o_data_a = 16'b1110001100001000;
            14'h29c1: o_data_a = 16'b0010100111000101;
            14'h29c2: o_data_a = 16'b1110110000010000;
            14'h29c3: o_data_a = 16'b0000000001011111;
            14'h29c4: o_data_a = 16'b1110101010000111;
            14'h29c5: o_data_a = 16'b0000000000000000;
            14'h29c6: o_data_a = 16'b1111110010101000;
            14'h29c7: o_data_a = 16'b1111110000010000;
            14'h29c8: o_data_a = 16'b0000000000000101;
            14'h29c9: o_data_a = 16'b1110001100001000;
            14'h29ca: o_data_a = 16'b0000000000101000;
            14'h29cb: o_data_a = 16'b1110110000010000;
            14'h29cc: o_data_a = 16'b0000000000000000;
            14'h29cd: o_data_a = 16'b1111110111101000;
            14'h29ce: o_data_a = 16'b1110110010100000;
            14'h29cf: o_data_a = 16'b1110001100001000;
            14'h29d0: o_data_a = 16'b0000000000011000;
            14'h29d1: o_data_a = 16'b1110110000010000;
            14'h29d2: o_data_a = 16'b0000000000000000;
            14'h29d3: o_data_a = 16'b1111110111101000;
            14'h29d4: o_data_a = 16'b1110110010100000;
            14'h29d5: o_data_a = 16'b1110001100001000;
            14'h29d6: o_data_a = 16'b0000000000001100;
            14'h29d7: o_data_a = 16'b1110110000010000;
            14'h29d8: o_data_a = 16'b0000000000000000;
            14'h29d9: o_data_a = 16'b1111110111101000;
            14'h29da: o_data_a = 16'b1110110010100000;
            14'h29db: o_data_a = 16'b1110001100001000;
            14'h29dc: o_data_a = 16'b0000000000000110;
            14'h29dd: o_data_a = 16'b1110110000010000;
            14'h29de: o_data_a = 16'b0000000000000000;
            14'h29df: o_data_a = 16'b1111110111101000;
            14'h29e0: o_data_a = 16'b1110110010100000;
            14'h29e1: o_data_a = 16'b1110001100001000;
            14'h29e2: o_data_a = 16'b0000000000000110;
            14'h29e3: o_data_a = 16'b1110110000010000;
            14'h29e4: o_data_a = 16'b0000000000000000;
            14'h29e5: o_data_a = 16'b1111110111101000;
            14'h29e6: o_data_a = 16'b1110110010100000;
            14'h29e7: o_data_a = 16'b1110001100001000;
            14'h29e8: o_data_a = 16'b0000000000000110;
            14'h29e9: o_data_a = 16'b1110110000010000;
            14'h29ea: o_data_a = 16'b0000000000000000;
            14'h29eb: o_data_a = 16'b1111110111101000;
            14'h29ec: o_data_a = 16'b1110110010100000;
            14'h29ed: o_data_a = 16'b1110001100001000;
            14'h29ee: o_data_a = 16'b0000000000000110;
            14'h29ef: o_data_a = 16'b1110110000010000;
            14'h29f0: o_data_a = 16'b0000000000000000;
            14'h29f1: o_data_a = 16'b1111110111101000;
            14'h29f2: o_data_a = 16'b1110110010100000;
            14'h29f3: o_data_a = 16'b1110001100001000;
            14'h29f4: o_data_a = 16'b0000000000000110;
            14'h29f5: o_data_a = 16'b1110110000010000;
            14'h29f6: o_data_a = 16'b0000000000000000;
            14'h29f7: o_data_a = 16'b1111110111101000;
            14'h29f8: o_data_a = 16'b1110110010100000;
            14'h29f9: o_data_a = 16'b1110001100001000;
            14'h29fa: o_data_a = 16'b0000000000001100;
            14'h29fb: o_data_a = 16'b1110110000010000;
            14'h29fc: o_data_a = 16'b0000000000000000;
            14'h29fd: o_data_a = 16'b1111110111101000;
            14'h29fe: o_data_a = 16'b1110110010100000;
            14'h29ff: o_data_a = 16'b1110001100001000;
            14'h2a00: o_data_a = 16'b0000000000011000;
            14'h2a01: o_data_a = 16'b1110110000010000;
            14'h2a02: o_data_a = 16'b0000000000000000;
            14'h2a03: o_data_a = 16'b1111110111101000;
            14'h2a04: o_data_a = 16'b1110110010100000;
            14'h2a05: o_data_a = 16'b1110001100001000;
            14'h2a06: o_data_a = 16'b0000000000000000;
            14'h2a07: o_data_a = 16'b1111110111001000;
            14'h2a08: o_data_a = 16'b1111110010100000;
            14'h2a09: o_data_a = 16'b1110101010001000;
            14'h2a0a: o_data_a = 16'b0000000000000000;
            14'h2a0b: o_data_a = 16'b1111110111001000;
            14'h2a0c: o_data_a = 16'b1111110010100000;
            14'h2a0d: o_data_a = 16'b1110101010001000;
            14'h2a0e: o_data_a = 16'b0000000000001100;
            14'h2a0f: o_data_a = 16'b1110110000010000;
            14'h2a10: o_data_a = 16'b0000000000001101;
            14'h2a11: o_data_a = 16'b1110001100001000;
            14'h2a12: o_data_a = 16'b0100010110110011;
            14'h2a13: o_data_a = 16'b1110110000010000;
            14'h2a14: o_data_a = 16'b0000000000001110;
            14'h2a15: o_data_a = 16'b1110001100001000;
            14'h2a16: o_data_a = 16'b0010101000011010;
            14'h2a17: o_data_a = 16'b1110110000010000;
            14'h2a18: o_data_a = 16'b0000000001011111;
            14'h2a19: o_data_a = 16'b1110101010000111;
            14'h2a1a: o_data_a = 16'b0000000000000000;
            14'h2a1b: o_data_a = 16'b1111110010101000;
            14'h2a1c: o_data_a = 16'b1111110000010000;
            14'h2a1d: o_data_a = 16'b0000000000000101;
            14'h2a1e: o_data_a = 16'b1110001100001000;
            14'h2a1f: o_data_a = 16'b0000000000101001;
            14'h2a20: o_data_a = 16'b1110110000010000;
            14'h2a21: o_data_a = 16'b0000000000000000;
            14'h2a22: o_data_a = 16'b1111110111101000;
            14'h2a23: o_data_a = 16'b1110110010100000;
            14'h2a24: o_data_a = 16'b1110001100001000;
            14'h2a25: o_data_a = 16'b0000000000000110;
            14'h2a26: o_data_a = 16'b1110110000010000;
            14'h2a27: o_data_a = 16'b0000000000000000;
            14'h2a28: o_data_a = 16'b1111110111101000;
            14'h2a29: o_data_a = 16'b1110110010100000;
            14'h2a2a: o_data_a = 16'b1110001100001000;
            14'h2a2b: o_data_a = 16'b0000000000001100;
            14'h2a2c: o_data_a = 16'b1110110000010000;
            14'h2a2d: o_data_a = 16'b0000000000000000;
            14'h2a2e: o_data_a = 16'b1111110111101000;
            14'h2a2f: o_data_a = 16'b1110110010100000;
            14'h2a30: o_data_a = 16'b1110001100001000;
            14'h2a31: o_data_a = 16'b0000000000011000;
            14'h2a32: o_data_a = 16'b1110110000010000;
            14'h2a33: o_data_a = 16'b0000000000000000;
            14'h2a34: o_data_a = 16'b1111110111101000;
            14'h2a35: o_data_a = 16'b1110110010100000;
            14'h2a36: o_data_a = 16'b1110001100001000;
            14'h2a37: o_data_a = 16'b0000000000011000;
            14'h2a38: o_data_a = 16'b1110110000010000;
            14'h2a39: o_data_a = 16'b0000000000000000;
            14'h2a3a: o_data_a = 16'b1111110111101000;
            14'h2a3b: o_data_a = 16'b1110110010100000;
            14'h2a3c: o_data_a = 16'b1110001100001000;
            14'h2a3d: o_data_a = 16'b0000000000011000;
            14'h2a3e: o_data_a = 16'b1110110000010000;
            14'h2a3f: o_data_a = 16'b0000000000000000;
            14'h2a40: o_data_a = 16'b1111110111101000;
            14'h2a41: o_data_a = 16'b1110110010100000;
            14'h2a42: o_data_a = 16'b1110001100001000;
            14'h2a43: o_data_a = 16'b0000000000011000;
            14'h2a44: o_data_a = 16'b1110110000010000;
            14'h2a45: o_data_a = 16'b0000000000000000;
            14'h2a46: o_data_a = 16'b1111110111101000;
            14'h2a47: o_data_a = 16'b1110110010100000;
            14'h2a48: o_data_a = 16'b1110001100001000;
            14'h2a49: o_data_a = 16'b0000000000011000;
            14'h2a4a: o_data_a = 16'b1110110000010000;
            14'h2a4b: o_data_a = 16'b0000000000000000;
            14'h2a4c: o_data_a = 16'b1111110111101000;
            14'h2a4d: o_data_a = 16'b1110110010100000;
            14'h2a4e: o_data_a = 16'b1110001100001000;
            14'h2a4f: o_data_a = 16'b0000000000001100;
            14'h2a50: o_data_a = 16'b1110110000010000;
            14'h2a51: o_data_a = 16'b0000000000000000;
            14'h2a52: o_data_a = 16'b1111110111101000;
            14'h2a53: o_data_a = 16'b1110110010100000;
            14'h2a54: o_data_a = 16'b1110001100001000;
            14'h2a55: o_data_a = 16'b0000000000000110;
            14'h2a56: o_data_a = 16'b1110110000010000;
            14'h2a57: o_data_a = 16'b0000000000000000;
            14'h2a58: o_data_a = 16'b1111110111101000;
            14'h2a59: o_data_a = 16'b1110110010100000;
            14'h2a5a: o_data_a = 16'b1110001100001000;
            14'h2a5b: o_data_a = 16'b0000000000000000;
            14'h2a5c: o_data_a = 16'b1111110111001000;
            14'h2a5d: o_data_a = 16'b1111110010100000;
            14'h2a5e: o_data_a = 16'b1110101010001000;
            14'h2a5f: o_data_a = 16'b0000000000000000;
            14'h2a60: o_data_a = 16'b1111110111001000;
            14'h2a61: o_data_a = 16'b1111110010100000;
            14'h2a62: o_data_a = 16'b1110101010001000;
            14'h2a63: o_data_a = 16'b0000000000001100;
            14'h2a64: o_data_a = 16'b1110110000010000;
            14'h2a65: o_data_a = 16'b0000000000001101;
            14'h2a66: o_data_a = 16'b1110001100001000;
            14'h2a67: o_data_a = 16'b0100010110110011;
            14'h2a68: o_data_a = 16'b1110110000010000;
            14'h2a69: o_data_a = 16'b0000000000001110;
            14'h2a6a: o_data_a = 16'b1110001100001000;
            14'h2a6b: o_data_a = 16'b0010101001101111;
            14'h2a6c: o_data_a = 16'b1110110000010000;
            14'h2a6d: o_data_a = 16'b0000000001011111;
            14'h2a6e: o_data_a = 16'b1110101010000111;
            14'h2a6f: o_data_a = 16'b0000000000000000;
            14'h2a70: o_data_a = 16'b1111110010101000;
            14'h2a71: o_data_a = 16'b1111110000010000;
            14'h2a72: o_data_a = 16'b0000000000000101;
            14'h2a73: o_data_a = 16'b1110001100001000;
            14'h2a74: o_data_a = 16'b0000000000101010;
            14'h2a75: o_data_a = 16'b1110110000010000;
            14'h2a76: o_data_a = 16'b0000000000000000;
            14'h2a77: o_data_a = 16'b1111110111101000;
            14'h2a78: o_data_a = 16'b1110110010100000;
            14'h2a79: o_data_a = 16'b1110001100001000;
            14'h2a7a: o_data_a = 16'b0000000000000000;
            14'h2a7b: o_data_a = 16'b1111110111001000;
            14'h2a7c: o_data_a = 16'b1111110010100000;
            14'h2a7d: o_data_a = 16'b1110101010001000;
            14'h2a7e: o_data_a = 16'b0000000000000000;
            14'h2a7f: o_data_a = 16'b1111110111001000;
            14'h2a80: o_data_a = 16'b1111110010100000;
            14'h2a81: o_data_a = 16'b1110101010001000;
            14'h2a82: o_data_a = 16'b0000000000000000;
            14'h2a83: o_data_a = 16'b1111110111001000;
            14'h2a84: o_data_a = 16'b1111110010100000;
            14'h2a85: o_data_a = 16'b1110101010001000;
            14'h2a86: o_data_a = 16'b0000000000110011;
            14'h2a87: o_data_a = 16'b1110110000010000;
            14'h2a88: o_data_a = 16'b0000000000000000;
            14'h2a89: o_data_a = 16'b1111110111101000;
            14'h2a8a: o_data_a = 16'b1110110010100000;
            14'h2a8b: o_data_a = 16'b1110001100001000;
            14'h2a8c: o_data_a = 16'b0000000000011110;
            14'h2a8d: o_data_a = 16'b1110110000010000;
            14'h2a8e: o_data_a = 16'b0000000000000000;
            14'h2a8f: o_data_a = 16'b1111110111101000;
            14'h2a90: o_data_a = 16'b1110110010100000;
            14'h2a91: o_data_a = 16'b1110001100001000;
            14'h2a92: o_data_a = 16'b0000000000111111;
            14'h2a93: o_data_a = 16'b1110110000010000;
            14'h2a94: o_data_a = 16'b0000000000000000;
            14'h2a95: o_data_a = 16'b1111110111101000;
            14'h2a96: o_data_a = 16'b1110110010100000;
            14'h2a97: o_data_a = 16'b1110001100001000;
            14'h2a98: o_data_a = 16'b0000000000011110;
            14'h2a99: o_data_a = 16'b1110110000010000;
            14'h2a9a: o_data_a = 16'b0000000000000000;
            14'h2a9b: o_data_a = 16'b1111110111101000;
            14'h2a9c: o_data_a = 16'b1110110010100000;
            14'h2a9d: o_data_a = 16'b1110001100001000;
            14'h2a9e: o_data_a = 16'b0000000000110011;
            14'h2a9f: o_data_a = 16'b1110110000010000;
            14'h2aa0: o_data_a = 16'b0000000000000000;
            14'h2aa1: o_data_a = 16'b1111110111101000;
            14'h2aa2: o_data_a = 16'b1110110010100000;
            14'h2aa3: o_data_a = 16'b1110001100001000;
            14'h2aa4: o_data_a = 16'b0000000000000000;
            14'h2aa5: o_data_a = 16'b1111110111001000;
            14'h2aa6: o_data_a = 16'b1111110010100000;
            14'h2aa7: o_data_a = 16'b1110101010001000;
            14'h2aa8: o_data_a = 16'b0000000000000000;
            14'h2aa9: o_data_a = 16'b1111110111001000;
            14'h2aaa: o_data_a = 16'b1111110010100000;
            14'h2aab: o_data_a = 16'b1110101010001000;
            14'h2aac: o_data_a = 16'b0000000000000000;
            14'h2aad: o_data_a = 16'b1111110111001000;
            14'h2aae: o_data_a = 16'b1111110010100000;
            14'h2aaf: o_data_a = 16'b1110101010001000;
            14'h2ab0: o_data_a = 16'b0000000000001100;
            14'h2ab1: o_data_a = 16'b1110110000010000;
            14'h2ab2: o_data_a = 16'b0000000000001101;
            14'h2ab3: o_data_a = 16'b1110001100001000;
            14'h2ab4: o_data_a = 16'b0100010110110011;
            14'h2ab5: o_data_a = 16'b1110110000010000;
            14'h2ab6: o_data_a = 16'b0000000000001110;
            14'h2ab7: o_data_a = 16'b1110001100001000;
            14'h2ab8: o_data_a = 16'b0010101010111100;
            14'h2ab9: o_data_a = 16'b1110110000010000;
            14'h2aba: o_data_a = 16'b0000000001011111;
            14'h2abb: o_data_a = 16'b1110101010000111;
            14'h2abc: o_data_a = 16'b0000000000000000;
            14'h2abd: o_data_a = 16'b1111110010101000;
            14'h2abe: o_data_a = 16'b1111110000010000;
            14'h2abf: o_data_a = 16'b0000000000000101;
            14'h2ac0: o_data_a = 16'b1110001100001000;
            14'h2ac1: o_data_a = 16'b0000000000101011;
            14'h2ac2: o_data_a = 16'b1110110000010000;
            14'h2ac3: o_data_a = 16'b0000000000000000;
            14'h2ac4: o_data_a = 16'b1111110111101000;
            14'h2ac5: o_data_a = 16'b1110110010100000;
            14'h2ac6: o_data_a = 16'b1110001100001000;
            14'h2ac7: o_data_a = 16'b0000000000000000;
            14'h2ac8: o_data_a = 16'b1111110111001000;
            14'h2ac9: o_data_a = 16'b1111110010100000;
            14'h2aca: o_data_a = 16'b1110101010001000;
            14'h2acb: o_data_a = 16'b0000000000000000;
            14'h2acc: o_data_a = 16'b1111110111001000;
            14'h2acd: o_data_a = 16'b1111110010100000;
            14'h2ace: o_data_a = 16'b1110101010001000;
            14'h2acf: o_data_a = 16'b0000000000000000;
            14'h2ad0: o_data_a = 16'b1111110111001000;
            14'h2ad1: o_data_a = 16'b1111110010100000;
            14'h2ad2: o_data_a = 16'b1110101010001000;
            14'h2ad3: o_data_a = 16'b0000000000001100;
            14'h2ad4: o_data_a = 16'b1110110000010000;
            14'h2ad5: o_data_a = 16'b0000000000000000;
            14'h2ad6: o_data_a = 16'b1111110111101000;
            14'h2ad7: o_data_a = 16'b1110110010100000;
            14'h2ad8: o_data_a = 16'b1110001100001000;
            14'h2ad9: o_data_a = 16'b0000000000001100;
            14'h2ada: o_data_a = 16'b1110110000010000;
            14'h2adb: o_data_a = 16'b0000000000000000;
            14'h2adc: o_data_a = 16'b1111110111101000;
            14'h2add: o_data_a = 16'b1110110010100000;
            14'h2ade: o_data_a = 16'b1110001100001000;
            14'h2adf: o_data_a = 16'b0000000000111111;
            14'h2ae0: o_data_a = 16'b1110110000010000;
            14'h2ae1: o_data_a = 16'b0000000000000000;
            14'h2ae2: o_data_a = 16'b1111110111101000;
            14'h2ae3: o_data_a = 16'b1110110010100000;
            14'h2ae4: o_data_a = 16'b1110001100001000;
            14'h2ae5: o_data_a = 16'b0000000000001100;
            14'h2ae6: o_data_a = 16'b1110110000010000;
            14'h2ae7: o_data_a = 16'b0000000000000000;
            14'h2ae8: o_data_a = 16'b1111110111101000;
            14'h2ae9: o_data_a = 16'b1110110010100000;
            14'h2aea: o_data_a = 16'b1110001100001000;
            14'h2aeb: o_data_a = 16'b0000000000001100;
            14'h2aec: o_data_a = 16'b1110110000010000;
            14'h2aed: o_data_a = 16'b0000000000000000;
            14'h2aee: o_data_a = 16'b1111110111101000;
            14'h2aef: o_data_a = 16'b1110110010100000;
            14'h2af0: o_data_a = 16'b1110001100001000;
            14'h2af1: o_data_a = 16'b0000000000000000;
            14'h2af2: o_data_a = 16'b1111110111001000;
            14'h2af3: o_data_a = 16'b1111110010100000;
            14'h2af4: o_data_a = 16'b1110101010001000;
            14'h2af5: o_data_a = 16'b0000000000000000;
            14'h2af6: o_data_a = 16'b1111110111001000;
            14'h2af7: o_data_a = 16'b1111110010100000;
            14'h2af8: o_data_a = 16'b1110101010001000;
            14'h2af9: o_data_a = 16'b0000000000000000;
            14'h2afa: o_data_a = 16'b1111110111001000;
            14'h2afb: o_data_a = 16'b1111110010100000;
            14'h2afc: o_data_a = 16'b1110101010001000;
            14'h2afd: o_data_a = 16'b0000000000001100;
            14'h2afe: o_data_a = 16'b1110110000010000;
            14'h2aff: o_data_a = 16'b0000000000001101;
            14'h2b00: o_data_a = 16'b1110001100001000;
            14'h2b01: o_data_a = 16'b0100010110110011;
            14'h2b02: o_data_a = 16'b1110110000010000;
            14'h2b03: o_data_a = 16'b0000000000001110;
            14'h2b04: o_data_a = 16'b1110001100001000;
            14'h2b05: o_data_a = 16'b0010101100001001;
            14'h2b06: o_data_a = 16'b1110110000010000;
            14'h2b07: o_data_a = 16'b0000000001011111;
            14'h2b08: o_data_a = 16'b1110101010000111;
            14'h2b09: o_data_a = 16'b0000000000000000;
            14'h2b0a: o_data_a = 16'b1111110010101000;
            14'h2b0b: o_data_a = 16'b1111110000010000;
            14'h2b0c: o_data_a = 16'b0000000000000101;
            14'h2b0d: o_data_a = 16'b1110001100001000;
            14'h2b0e: o_data_a = 16'b0000000000101100;
            14'h2b0f: o_data_a = 16'b1110110000010000;
            14'h2b10: o_data_a = 16'b0000000000000000;
            14'h2b11: o_data_a = 16'b1111110111101000;
            14'h2b12: o_data_a = 16'b1110110010100000;
            14'h2b13: o_data_a = 16'b1110001100001000;
            14'h2b14: o_data_a = 16'b0000000000000000;
            14'h2b15: o_data_a = 16'b1111110111001000;
            14'h2b16: o_data_a = 16'b1111110010100000;
            14'h2b17: o_data_a = 16'b1110101010001000;
            14'h2b18: o_data_a = 16'b0000000000000000;
            14'h2b19: o_data_a = 16'b1111110111001000;
            14'h2b1a: o_data_a = 16'b1111110010100000;
            14'h2b1b: o_data_a = 16'b1110101010001000;
            14'h2b1c: o_data_a = 16'b0000000000000000;
            14'h2b1d: o_data_a = 16'b1111110111001000;
            14'h2b1e: o_data_a = 16'b1111110010100000;
            14'h2b1f: o_data_a = 16'b1110101010001000;
            14'h2b20: o_data_a = 16'b0000000000000000;
            14'h2b21: o_data_a = 16'b1111110111001000;
            14'h2b22: o_data_a = 16'b1111110010100000;
            14'h2b23: o_data_a = 16'b1110101010001000;
            14'h2b24: o_data_a = 16'b0000000000000000;
            14'h2b25: o_data_a = 16'b1111110111001000;
            14'h2b26: o_data_a = 16'b1111110010100000;
            14'h2b27: o_data_a = 16'b1110101010001000;
            14'h2b28: o_data_a = 16'b0000000000000000;
            14'h2b29: o_data_a = 16'b1111110111001000;
            14'h2b2a: o_data_a = 16'b1111110010100000;
            14'h2b2b: o_data_a = 16'b1110101010001000;
            14'h2b2c: o_data_a = 16'b0000000000000000;
            14'h2b2d: o_data_a = 16'b1111110111001000;
            14'h2b2e: o_data_a = 16'b1111110010100000;
            14'h2b2f: o_data_a = 16'b1110101010001000;
            14'h2b30: o_data_a = 16'b0000000000001100;
            14'h2b31: o_data_a = 16'b1110110000010000;
            14'h2b32: o_data_a = 16'b0000000000000000;
            14'h2b33: o_data_a = 16'b1111110111101000;
            14'h2b34: o_data_a = 16'b1110110010100000;
            14'h2b35: o_data_a = 16'b1110001100001000;
            14'h2b36: o_data_a = 16'b0000000000001100;
            14'h2b37: o_data_a = 16'b1110110000010000;
            14'h2b38: o_data_a = 16'b0000000000000000;
            14'h2b39: o_data_a = 16'b1111110111101000;
            14'h2b3a: o_data_a = 16'b1110110010100000;
            14'h2b3b: o_data_a = 16'b1110001100001000;
            14'h2b3c: o_data_a = 16'b0000000000000110;
            14'h2b3d: o_data_a = 16'b1110110000010000;
            14'h2b3e: o_data_a = 16'b0000000000000000;
            14'h2b3f: o_data_a = 16'b1111110111101000;
            14'h2b40: o_data_a = 16'b1110110010100000;
            14'h2b41: o_data_a = 16'b1110001100001000;
            14'h2b42: o_data_a = 16'b0000000000000000;
            14'h2b43: o_data_a = 16'b1111110111001000;
            14'h2b44: o_data_a = 16'b1111110010100000;
            14'h2b45: o_data_a = 16'b1110101010001000;
            14'h2b46: o_data_a = 16'b0000000000001100;
            14'h2b47: o_data_a = 16'b1110110000010000;
            14'h2b48: o_data_a = 16'b0000000000001101;
            14'h2b49: o_data_a = 16'b1110001100001000;
            14'h2b4a: o_data_a = 16'b0100010110110011;
            14'h2b4b: o_data_a = 16'b1110110000010000;
            14'h2b4c: o_data_a = 16'b0000000000001110;
            14'h2b4d: o_data_a = 16'b1110001100001000;
            14'h2b4e: o_data_a = 16'b0010101101010010;
            14'h2b4f: o_data_a = 16'b1110110000010000;
            14'h2b50: o_data_a = 16'b0000000001011111;
            14'h2b51: o_data_a = 16'b1110101010000111;
            14'h2b52: o_data_a = 16'b0000000000000000;
            14'h2b53: o_data_a = 16'b1111110010101000;
            14'h2b54: o_data_a = 16'b1111110000010000;
            14'h2b55: o_data_a = 16'b0000000000000101;
            14'h2b56: o_data_a = 16'b1110001100001000;
            14'h2b57: o_data_a = 16'b0000000000101101;
            14'h2b58: o_data_a = 16'b1110110000010000;
            14'h2b59: o_data_a = 16'b0000000000000000;
            14'h2b5a: o_data_a = 16'b1111110111101000;
            14'h2b5b: o_data_a = 16'b1110110010100000;
            14'h2b5c: o_data_a = 16'b1110001100001000;
            14'h2b5d: o_data_a = 16'b0000000000000000;
            14'h2b5e: o_data_a = 16'b1111110111001000;
            14'h2b5f: o_data_a = 16'b1111110010100000;
            14'h2b60: o_data_a = 16'b1110101010001000;
            14'h2b61: o_data_a = 16'b0000000000000000;
            14'h2b62: o_data_a = 16'b1111110111001000;
            14'h2b63: o_data_a = 16'b1111110010100000;
            14'h2b64: o_data_a = 16'b1110101010001000;
            14'h2b65: o_data_a = 16'b0000000000000000;
            14'h2b66: o_data_a = 16'b1111110111001000;
            14'h2b67: o_data_a = 16'b1111110010100000;
            14'h2b68: o_data_a = 16'b1110101010001000;
            14'h2b69: o_data_a = 16'b0000000000000000;
            14'h2b6a: o_data_a = 16'b1111110111001000;
            14'h2b6b: o_data_a = 16'b1111110010100000;
            14'h2b6c: o_data_a = 16'b1110101010001000;
            14'h2b6d: o_data_a = 16'b0000000000000000;
            14'h2b6e: o_data_a = 16'b1111110111001000;
            14'h2b6f: o_data_a = 16'b1111110010100000;
            14'h2b70: o_data_a = 16'b1110101010001000;
            14'h2b71: o_data_a = 16'b0000000000111111;
            14'h2b72: o_data_a = 16'b1110110000010000;
            14'h2b73: o_data_a = 16'b0000000000000000;
            14'h2b74: o_data_a = 16'b1111110111101000;
            14'h2b75: o_data_a = 16'b1110110010100000;
            14'h2b76: o_data_a = 16'b1110001100001000;
            14'h2b77: o_data_a = 16'b0000000000000000;
            14'h2b78: o_data_a = 16'b1111110111001000;
            14'h2b79: o_data_a = 16'b1111110010100000;
            14'h2b7a: o_data_a = 16'b1110101010001000;
            14'h2b7b: o_data_a = 16'b0000000000000000;
            14'h2b7c: o_data_a = 16'b1111110111001000;
            14'h2b7d: o_data_a = 16'b1111110010100000;
            14'h2b7e: o_data_a = 16'b1110101010001000;
            14'h2b7f: o_data_a = 16'b0000000000000000;
            14'h2b80: o_data_a = 16'b1111110111001000;
            14'h2b81: o_data_a = 16'b1111110010100000;
            14'h2b82: o_data_a = 16'b1110101010001000;
            14'h2b83: o_data_a = 16'b0000000000000000;
            14'h2b84: o_data_a = 16'b1111110111001000;
            14'h2b85: o_data_a = 16'b1111110010100000;
            14'h2b86: o_data_a = 16'b1110101010001000;
            14'h2b87: o_data_a = 16'b0000000000000000;
            14'h2b88: o_data_a = 16'b1111110111001000;
            14'h2b89: o_data_a = 16'b1111110010100000;
            14'h2b8a: o_data_a = 16'b1110101010001000;
            14'h2b8b: o_data_a = 16'b0000000000001100;
            14'h2b8c: o_data_a = 16'b1110110000010000;
            14'h2b8d: o_data_a = 16'b0000000000001101;
            14'h2b8e: o_data_a = 16'b1110001100001000;
            14'h2b8f: o_data_a = 16'b0100010110110011;
            14'h2b90: o_data_a = 16'b1110110000010000;
            14'h2b91: o_data_a = 16'b0000000000001110;
            14'h2b92: o_data_a = 16'b1110001100001000;
            14'h2b93: o_data_a = 16'b0010101110010111;
            14'h2b94: o_data_a = 16'b1110110000010000;
            14'h2b95: o_data_a = 16'b0000000001011111;
            14'h2b96: o_data_a = 16'b1110101010000111;
            14'h2b97: o_data_a = 16'b0000000000000000;
            14'h2b98: o_data_a = 16'b1111110010101000;
            14'h2b99: o_data_a = 16'b1111110000010000;
            14'h2b9a: o_data_a = 16'b0000000000000101;
            14'h2b9b: o_data_a = 16'b1110001100001000;
            14'h2b9c: o_data_a = 16'b0000000000101110;
            14'h2b9d: o_data_a = 16'b1110110000010000;
            14'h2b9e: o_data_a = 16'b0000000000000000;
            14'h2b9f: o_data_a = 16'b1111110111101000;
            14'h2ba0: o_data_a = 16'b1110110010100000;
            14'h2ba1: o_data_a = 16'b1110001100001000;
            14'h2ba2: o_data_a = 16'b0000000000000000;
            14'h2ba3: o_data_a = 16'b1111110111001000;
            14'h2ba4: o_data_a = 16'b1111110010100000;
            14'h2ba5: o_data_a = 16'b1110101010001000;
            14'h2ba6: o_data_a = 16'b0000000000000000;
            14'h2ba7: o_data_a = 16'b1111110111001000;
            14'h2ba8: o_data_a = 16'b1111110010100000;
            14'h2ba9: o_data_a = 16'b1110101010001000;
            14'h2baa: o_data_a = 16'b0000000000000000;
            14'h2bab: o_data_a = 16'b1111110111001000;
            14'h2bac: o_data_a = 16'b1111110010100000;
            14'h2bad: o_data_a = 16'b1110101010001000;
            14'h2bae: o_data_a = 16'b0000000000000000;
            14'h2baf: o_data_a = 16'b1111110111001000;
            14'h2bb0: o_data_a = 16'b1111110010100000;
            14'h2bb1: o_data_a = 16'b1110101010001000;
            14'h2bb2: o_data_a = 16'b0000000000000000;
            14'h2bb3: o_data_a = 16'b1111110111001000;
            14'h2bb4: o_data_a = 16'b1111110010100000;
            14'h2bb5: o_data_a = 16'b1110101010001000;
            14'h2bb6: o_data_a = 16'b0000000000000000;
            14'h2bb7: o_data_a = 16'b1111110111001000;
            14'h2bb8: o_data_a = 16'b1111110010100000;
            14'h2bb9: o_data_a = 16'b1110101010001000;
            14'h2bba: o_data_a = 16'b0000000000000000;
            14'h2bbb: o_data_a = 16'b1111110111001000;
            14'h2bbc: o_data_a = 16'b1111110010100000;
            14'h2bbd: o_data_a = 16'b1110101010001000;
            14'h2bbe: o_data_a = 16'b0000000000001100;
            14'h2bbf: o_data_a = 16'b1110110000010000;
            14'h2bc0: o_data_a = 16'b0000000000000000;
            14'h2bc1: o_data_a = 16'b1111110111101000;
            14'h2bc2: o_data_a = 16'b1110110010100000;
            14'h2bc3: o_data_a = 16'b1110001100001000;
            14'h2bc4: o_data_a = 16'b0000000000001100;
            14'h2bc5: o_data_a = 16'b1110110000010000;
            14'h2bc6: o_data_a = 16'b0000000000000000;
            14'h2bc7: o_data_a = 16'b1111110111101000;
            14'h2bc8: o_data_a = 16'b1110110010100000;
            14'h2bc9: o_data_a = 16'b1110001100001000;
            14'h2bca: o_data_a = 16'b0000000000000000;
            14'h2bcb: o_data_a = 16'b1111110111001000;
            14'h2bcc: o_data_a = 16'b1111110010100000;
            14'h2bcd: o_data_a = 16'b1110101010001000;
            14'h2bce: o_data_a = 16'b0000000000000000;
            14'h2bcf: o_data_a = 16'b1111110111001000;
            14'h2bd0: o_data_a = 16'b1111110010100000;
            14'h2bd1: o_data_a = 16'b1110101010001000;
            14'h2bd2: o_data_a = 16'b0000000000001100;
            14'h2bd3: o_data_a = 16'b1110110000010000;
            14'h2bd4: o_data_a = 16'b0000000000001101;
            14'h2bd5: o_data_a = 16'b1110001100001000;
            14'h2bd6: o_data_a = 16'b0100010110110011;
            14'h2bd7: o_data_a = 16'b1110110000010000;
            14'h2bd8: o_data_a = 16'b0000000000001110;
            14'h2bd9: o_data_a = 16'b1110001100001000;
            14'h2bda: o_data_a = 16'b0010101111011110;
            14'h2bdb: o_data_a = 16'b1110110000010000;
            14'h2bdc: o_data_a = 16'b0000000001011111;
            14'h2bdd: o_data_a = 16'b1110101010000111;
            14'h2bde: o_data_a = 16'b0000000000000000;
            14'h2bdf: o_data_a = 16'b1111110010101000;
            14'h2be0: o_data_a = 16'b1111110000010000;
            14'h2be1: o_data_a = 16'b0000000000000101;
            14'h2be2: o_data_a = 16'b1110001100001000;
            14'h2be3: o_data_a = 16'b0000000000101111;
            14'h2be4: o_data_a = 16'b1110110000010000;
            14'h2be5: o_data_a = 16'b0000000000000000;
            14'h2be6: o_data_a = 16'b1111110111101000;
            14'h2be7: o_data_a = 16'b1110110010100000;
            14'h2be8: o_data_a = 16'b1110001100001000;
            14'h2be9: o_data_a = 16'b0000000000000000;
            14'h2bea: o_data_a = 16'b1111110111001000;
            14'h2beb: o_data_a = 16'b1111110010100000;
            14'h2bec: o_data_a = 16'b1110101010001000;
            14'h2bed: o_data_a = 16'b0000000000000000;
            14'h2bee: o_data_a = 16'b1111110111001000;
            14'h2bef: o_data_a = 16'b1111110010100000;
            14'h2bf0: o_data_a = 16'b1110101010001000;
            14'h2bf1: o_data_a = 16'b0000000000100000;
            14'h2bf2: o_data_a = 16'b1110110000010000;
            14'h2bf3: o_data_a = 16'b0000000000000000;
            14'h2bf4: o_data_a = 16'b1111110111101000;
            14'h2bf5: o_data_a = 16'b1110110010100000;
            14'h2bf6: o_data_a = 16'b1110001100001000;
            14'h2bf7: o_data_a = 16'b0000000000110000;
            14'h2bf8: o_data_a = 16'b1110110000010000;
            14'h2bf9: o_data_a = 16'b0000000000000000;
            14'h2bfa: o_data_a = 16'b1111110111101000;
            14'h2bfb: o_data_a = 16'b1110110010100000;
            14'h2bfc: o_data_a = 16'b1110001100001000;
            14'h2bfd: o_data_a = 16'b0000000000011000;
            14'h2bfe: o_data_a = 16'b1110110000010000;
            14'h2bff: o_data_a = 16'b0000000000000000;
            14'h2c00: o_data_a = 16'b1111110111101000;
            14'h2c01: o_data_a = 16'b1110110010100000;
            14'h2c02: o_data_a = 16'b1110001100001000;
            14'h2c03: o_data_a = 16'b0000000000001100;
            14'h2c04: o_data_a = 16'b1110110000010000;
            14'h2c05: o_data_a = 16'b0000000000000000;
            14'h2c06: o_data_a = 16'b1111110111101000;
            14'h2c07: o_data_a = 16'b1110110010100000;
            14'h2c08: o_data_a = 16'b1110001100001000;
            14'h2c09: o_data_a = 16'b0000000000000110;
            14'h2c0a: o_data_a = 16'b1110110000010000;
            14'h2c0b: o_data_a = 16'b0000000000000000;
            14'h2c0c: o_data_a = 16'b1111110111101000;
            14'h2c0d: o_data_a = 16'b1110110010100000;
            14'h2c0e: o_data_a = 16'b1110001100001000;
            14'h2c0f: o_data_a = 16'b0000000000000011;
            14'h2c10: o_data_a = 16'b1110110000010000;
            14'h2c11: o_data_a = 16'b0000000000000000;
            14'h2c12: o_data_a = 16'b1111110111101000;
            14'h2c13: o_data_a = 16'b1110110010100000;
            14'h2c14: o_data_a = 16'b1110001100001000;
            14'h2c15: o_data_a = 16'b0000000000000000;
            14'h2c16: o_data_a = 16'b1111110111001000;
            14'h2c17: o_data_a = 16'b1111110010100000;
            14'h2c18: o_data_a = 16'b1110111111001000;
            14'h2c19: o_data_a = 16'b0000000000000000;
            14'h2c1a: o_data_a = 16'b1111110111001000;
            14'h2c1b: o_data_a = 16'b1111110010100000;
            14'h2c1c: o_data_a = 16'b1110101010001000;
            14'h2c1d: o_data_a = 16'b0000000000000000;
            14'h2c1e: o_data_a = 16'b1111110111001000;
            14'h2c1f: o_data_a = 16'b1111110010100000;
            14'h2c20: o_data_a = 16'b1110101010001000;
            14'h2c21: o_data_a = 16'b0000000000001100;
            14'h2c22: o_data_a = 16'b1110110000010000;
            14'h2c23: o_data_a = 16'b0000000000001101;
            14'h2c24: o_data_a = 16'b1110001100001000;
            14'h2c25: o_data_a = 16'b0100010110110011;
            14'h2c26: o_data_a = 16'b1110110000010000;
            14'h2c27: o_data_a = 16'b0000000000001110;
            14'h2c28: o_data_a = 16'b1110001100001000;
            14'h2c29: o_data_a = 16'b0010110000101101;
            14'h2c2a: o_data_a = 16'b1110110000010000;
            14'h2c2b: o_data_a = 16'b0000000001011111;
            14'h2c2c: o_data_a = 16'b1110101010000111;
            14'h2c2d: o_data_a = 16'b0000000000000000;
            14'h2c2e: o_data_a = 16'b1111110010101000;
            14'h2c2f: o_data_a = 16'b1111110000010000;
            14'h2c30: o_data_a = 16'b0000000000000101;
            14'h2c31: o_data_a = 16'b1110001100001000;
            14'h2c32: o_data_a = 16'b0000000000110000;
            14'h2c33: o_data_a = 16'b1110110000010000;
            14'h2c34: o_data_a = 16'b0000000000000000;
            14'h2c35: o_data_a = 16'b1111110111101000;
            14'h2c36: o_data_a = 16'b1110110010100000;
            14'h2c37: o_data_a = 16'b1110001100001000;
            14'h2c38: o_data_a = 16'b0000000000001100;
            14'h2c39: o_data_a = 16'b1110110000010000;
            14'h2c3a: o_data_a = 16'b0000000000000000;
            14'h2c3b: o_data_a = 16'b1111110111101000;
            14'h2c3c: o_data_a = 16'b1110110010100000;
            14'h2c3d: o_data_a = 16'b1110001100001000;
            14'h2c3e: o_data_a = 16'b0000000000011110;
            14'h2c3f: o_data_a = 16'b1110110000010000;
            14'h2c40: o_data_a = 16'b0000000000000000;
            14'h2c41: o_data_a = 16'b1111110111101000;
            14'h2c42: o_data_a = 16'b1110110010100000;
            14'h2c43: o_data_a = 16'b1110001100001000;
            14'h2c44: o_data_a = 16'b0000000000110011;
            14'h2c45: o_data_a = 16'b1110110000010000;
            14'h2c46: o_data_a = 16'b0000000000000000;
            14'h2c47: o_data_a = 16'b1111110111101000;
            14'h2c48: o_data_a = 16'b1110110010100000;
            14'h2c49: o_data_a = 16'b1110001100001000;
            14'h2c4a: o_data_a = 16'b0000000000110011;
            14'h2c4b: o_data_a = 16'b1110110000010000;
            14'h2c4c: o_data_a = 16'b0000000000000000;
            14'h2c4d: o_data_a = 16'b1111110111101000;
            14'h2c4e: o_data_a = 16'b1110110010100000;
            14'h2c4f: o_data_a = 16'b1110001100001000;
            14'h2c50: o_data_a = 16'b0000000000110011;
            14'h2c51: o_data_a = 16'b1110110000010000;
            14'h2c52: o_data_a = 16'b0000000000000000;
            14'h2c53: o_data_a = 16'b1111110111101000;
            14'h2c54: o_data_a = 16'b1110110010100000;
            14'h2c55: o_data_a = 16'b1110001100001000;
            14'h2c56: o_data_a = 16'b0000000000110011;
            14'h2c57: o_data_a = 16'b1110110000010000;
            14'h2c58: o_data_a = 16'b0000000000000000;
            14'h2c59: o_data_a = 16'b1111110111101000;
            14'h2c5a: o_data_a = 16'b1110110010100000;
            14'h2c5b: o_data_a = 16'b1110001100001000;
            14'h2c5c: o_data_a = 16'b0000000000110011;
            14'h2c5d: o_data_a = 16'b1110110000010000;
            14'h2c5e: o_data_a = 16'b0000000000000000;
            14'h2c5f: o_data_a = 16'b1111110111101000;
            14'h2c60: o_data_a = 16'b1110110010100000;
            14'h2c61: o_data_a = 16'b1110001100001000;
            14'h2c62: o_data_a = 16'b0000000000011110;
            14'h2c63: o_data_a = 16'b1110110000010000;
            14'h2c64: o_data_a = 16'b0000000000000000;
            14'h2c65: o_data_a = 16'b1111110111101000;
            14'h2c66: o_data_a = 16'b1110110010100000;
            14'h2c67: o_data_a = 16'b1110001100001000;
            14'h2c68: o_data_a = 16'b0000000000001100;
            14'h2c69: o_data_a = 16'b1110110000010000;
            14'h2c6a: o_data_a = 16'b0000000000000000;
            14'h2c6b: o_data_a = 16'b1111110111101000;
            14'h2c6c: o_data_a = 16'b1110110010100000;
            14'h2c6d: o_data_a = 16'b1110001100001000;
            14'h2c6e: o_data_a = 16'b0000000000000000;
            14'h2c6f: o_data_a = 16'b1111110111001000;
            14'h2c70: o_data_a = 16'b1111110010100000;
            14'h2c71: o_data_a = 16'b1110101010001000;
            14'h2c72: o_data_a = 16'b0000000000000000;
            14'h2c73: o_data_a = 16'b1111110111001000;
            14'h2c74: o_data_a = 16'b1111110010100000;
            14'h2c75: o_data_a = 16'b1110101010001000;
            14'h2c76: o_data_a = 16'b0000000000001100;
            14'h2c77: o_data_a = 16'b1110110000010000;
            14'h2c78: o_data_a = 16'b0000000000001101;
            14'h2c79: o_data_a = 16'b1110001100001000;
            14'h2c7a: o_data_a = 16'b0100010110110011;
            14'h2c7b: o_data_a = 16'b1110110000010000;
            14'h2c7c: o_data_a = 16'b0000000000001110;
            14'h2c7d: o_data_a = 16'b1110001100001000;
            14'h2c7e: o_data_a = 16'b0010110010000010;
            14'h2c7f: o_data_a = 16'b1110110000010000;
            14'h2c80: o_data_a = 16'b0000000001011111;
            14'h2c81: o_data_a = 16'b1110101010000111;
            14'h2c82: o_data_a = 16'b0000000000000000;
            14'h2c83: o_data_a = 16'b1111110010101000;
            14'h2c84: o_data_a = 16'b1111110000010000;
            14'h2c85: o_data_a = 16'b0000000000000101;
            14'h2c86: o_data_a = 16'b1110001100001000;
            14'h2c87: o_data_a = 16'b0000000000110001;
            14'h2c88: o_data_a = 16'b1110110000010000;
            14'h2c89: o_data_a = 16'b0000000000000000;
            14'h2c8a: o_data_a = 16'b1111110111101000;
            14'h2c8b: o_data_a = 16'b1110110010100000;
            14'h2c8c: o_data_a = 16'b1110001100001000;
            14'h2c8d: o_data_a = 16'b0000000000001100;
            14'h2c8e: o_data_a = 16'b1110110000010000;
            14'h2c8f: o_data_a = 16'b0000000000000000;
            14'h2c90: o_data_a = 16'b1111110111101000;
            14'h2c91: o_data_a = 16'b1110110010100000;
            14'h2c92: o_data_a = 16'b1110001100001000;
            14'h2c93: o_data_a = 16'b0000000000001110;
            14'h2c94: o_data_a = 16'b1110110000010000;
            14'h2c95: o_data_a = 16'b0000000000000000;
            14'h2c96: o_data_a = 16'b1111110111101000;
            14'h2c97: o_data_a = 16'b1110110010100000;
            14'h2c98: o_data_a = 16'b1110001100001000;
            14'h2c99: o_data_a = 16'b0000000000001111;
            14'h2c9a: o_data_a = 16'b1110110000010000;
            14'h2c9b: o_data_a = 16'b0000000000000000;
            14'h2c9c: o_data_a = 16'b1111110111101000;
            14'h2c9d: o_data_a = 16'b1110110010100000;
            14'h2c9e: o_data_a = 16'b1110001100001000;
            14'h2c9f: o_data_a = 16'b0000000000001100;
            14'h2ca0: o_data_a = 16'b1110110000010000;
            14'h2ca1: o_data_a = 16'b0000000000000000;
            14'h2ca2: o_data_a = 16'b1111110111101000;
            14'h2ca3: o_data_a = 16'b1110110010100000;
            14'h2ca4: o_data_a = 16'b1110001100001000;
            14'h2ca5: o_data_a = 16'b0000000000001100;
            14'h2ca6: o_data_a = 16'b1110110000010000;
            14'h2ca7: o_data_a = 16'b0000000000000000;
            14'h2ca8: o_data_a = 16'b1111110111101000;
            14'h2ca9: o_data_a = 16'b1110110010100000;
            14'h2caa: o_data_a = 16'b1110001100001000;
            14'h2cab: o_data_a = 16'b0000000000001100;
            14'h2cac: o_data_a = 16'b1110110000010000;
            14'h2cad: o_data_a = 16'b0000000000000000;
            14'h2cae: o_data_a = 16'b1111110111101000;
            14'h2caf: o_data_a = 16'b1110110010100000;
            14'h2cb0: o_data_a = 16'b1110001100001000;
            14'h2cb1: o_data_a = 16'b0000000000001100;
            14'h2cb2: o_data_a = 16'b1110110000010000;
            14'h2cb3: o_data_a = 16'b0000000000000000;
            14'h2cb4: o_data_a = 16'b1111110111101000;
            14'h2cb5: o_data_a = 16'b1110110010100000;
            14'h2cb6: o_data_a = 16'b1110001100001000;
            14'h2cb7: o_data_a = 16'b0000000000001100;
            14'h2cb8: o_data_a = 16'b1110110000010000;
            14'h2cb9: o_data_a = 16'b0000000000000000;
            14'h2cba: o_data_a = 16'b1111110111101000;
            14'h2cbb: o_data_a = 16'b1110110010100000;
            14'h2cbc: o_data_a = 16'b1110001100001000;
            14'h2cbd: o_data_a = 16'b0000000000111111;
            14'h2cbe: o_data_a = 16'b1110110000010000;
            14'h2cbf: o_data_a = 16'b0000000000000000;
            14'h2cc0: o_data_a = 16'b1111110111101000;
            14'h2cc1: o_data_a = 16'b1110110010100000;
            14'h2cc2: o_data_a = 16'b1110001100001000;
            14'h2cc3: o_data_a = 16'b0000000000000000;
            14'h2cc4: o_data_a = 16'b1111110111001000;
            14'h2cc5: o_data_a = 16'b1111110010100000;
            14'h2cc6: o_data_a = 16'b1110101010001000;
            14'h2cc7: o_data_a = 16'b0000000000000000;
            14'h2cc8: o_data_a = 16'b1111110111001000;
            14'h2cc9: o_data_a = 16'b1111110010100000;
            14'h2cca: o_data_a = 16'b1110101010001000;
            14'h2ccb: o_data_a = 16'b0000000000001100;
            14'h2ccc: o_data_a = 16'b1110110000010000;
            14'h2ccd: o_data_a = 16'b0000000000001101;
            14'h2cce: o_data_a = 16'b1110001100001000;
            14'h2ccf: o_data_a = 16'b0100010110110011;
            14'h2cd0: o_data_a = 16'b1110110000010000;
            14'h2cd1: o_data_a = 16'b0000000000001110;
            14'h2cd2: o_data_a = 16'b1110001100001000;
            14'h2cd3: o_data_a = 16'b0010110011010111;
            14'h2cd4: o_data_a = 16'b1110110000010000;
            14'h2cd5: o_data_a = 16'b0000000001011111;
            14'h2cd6: o_data_a = 16'b1110101010000111;
            14'h2cd7: o_data_a = 16'b0000000000000000;
            14'h2cd8: o_data_a = 16'b1111110010101000;
            14'h2cd9: o_data_a = 16'b1111110000010000;
            14'h2cda: o_data_a = 16'b0000000000000101;
            14'h2cdb: o_data_a = 16'b1110001100001000;
            14'h2cdc: o_data_a = 16'b0000000000110010;
            14'h2cdd: o_data_a = 16'b1110110000010000;
            14'h2cde: o_data_a = 16'b0000000000000000;
            14'h2cdf: o_data_a = 16'b1111110111101000;
            14'h2ce0: o_data_a = 16'b1110110010100000;
            14'h2ce1: o_data_a = 16'b1110001100001000;
            14'h2ce2: o_data_a = 16'b0000000000011110;
            14'h2ce3: o_data_a = 16'b1110110000010000;
            14'h2ce4: o_data_a = 16'b0000000000000000;
            14'h2ce5: o_data_a = 16'b1111110111101000;
            14'h2ce6: o_data_a = 16'b1110110010100000;
            14'h2ce7: o_data_a = 16'b1110001100001000;
            14'h2ce8: o_data_a = 16'b0000000000110011;
            14'h2ce9: o_data_a = 16'b1110110000010000;
            14'h2cea: o_data_a = 16'b0000000000000000;
            14'h2ceb: o_data_a = 16'b1111110111101000;
            14'h2cec: o_data_a = 16'b1110110010100000;
            14'h2ced: o_data_a = 16'b1110001100001000;
            14'h2cee: o_data_a = 16'b0000000000110000;
            14'h2cef: o_data_a = 16'b1110110000010000;
            14'h2cf0: o_data_a = 16'b0000000000000000;
            14'h2cf1: o_data_a = 16'b1111110111101000;
            14'h2cf2: o_data_a = 16'b1110110010100000;
            14'h2cf3: o_data_a = 16'b1110001100001000;
            14'h2cf4: o_data_a = 16'b0000000000011000;
            14'h2cf5: o_data_a = 16'b1110110000010000;
            14'h2cf6: o_data_a = 16'b0000000000000000;
            14'h2cf7: o_data_a = 16'b1111110111101000;
            14'h2cf8: o_data_a = 16'b1110110010100000;
            14'h2cf9: o_data_a = 16'b1110001100001000;
            14'h2cfa: o_data_a = 16'b0000000000001100;
            14'h2cfb: o_data_a = 16'b1110110000010000;
            14'h2cfc: o_data_a = 16'b0000000000000000;
            14'h2cfd: o_data_a = 16'b1111110111101000;
            14'h2cfe: o_data_a = 16'b1110110010100000;
            14'h2cff: o_data_a = 16'b1110001100001000;
            14'h2d00: o_data_a = 16'b0000000000000110;
            14'h2d01: o_data_a = 16'b1110110000010000;
            14'h2d02: o_data_a = 16'b0000000000000000;
            14'h2d03: o_data_a = 16'b1111110111101000;
            14'h2d04: o_data_a = 16'b1110110010100000;
            14'h2d05: o_data_a = 16'b1110001100001000;
            14'h2d06: o_data_a = 16'b0000000000000011;
            14'h2d07: o_data_a = 16'b1110110000010000;
            14'h2d08: o_data_a = 16'b0000000000000000;
            14'h2d09: o_data_a = 16'b1111110111101000;
            14'h2d0a: o_data_a = 16'b1110110010100000;
            14'h2d0b: o_data_a = 16'b1110001100001000;
            14'h2d0c: o_data_a = 16'b0000000000110011;
            14'h2d0d: o_data_a = 16'b1110110000010000;
            14'h2d0e: o_data_a = 16'b0000000000000000;
            14'h2d0f: o_data_a = 16'b1111110111101000;
            14'h2d10: o_data_a = 16'b1110110010100000;
            14'h2d11: o_data_a = 16'b1110001100001000;
            14'h2d12: o_data_a = 16'b0000000000111111;
            14'h2d13: o_data_a = 16'b1110110000010000;
            14'h2d14: o_data_a = 16'b0000000000000000;
            14'h2d15: o_data_a = 16'b1111110111101000;
            14'h2d16: o_data_a = 16'b1110110010100000;
            14'h2d17: o_data_a = 16'b1110001100001000;
            14'h2d18: o_data_a = 16'b0000000000000000;
            14'h2d19: o_data_a = 16'b1111110111001000;
            14'h2d1a: o_data_a = 16'b1111110010100000;
            14'h2d1b: o_data_a = 16'b1110101010001000;
            14'h2d1c: o_data_a = 16'b0000000000000000;
            14'h2d1d: o_data_a = 16'b1111110111001000;
            14'h2d1e: o_data_a = 16'b1111110010100000;
            14'h2d1f: o_data_a = 16'b1110101010001000;
            14'h2d20: o_data_a = 16'b0000000000001100;
            14'h2d21: o_data_a = 16'b1110110000010000;
            14'h2d22: o_data_a = 16'b0000000000001101;
            14'h2d23: o_data_a = 16'b1110001100001000;
            14'h2d24: o_data_a = 16'b0100010110110011;
            14'h2d25: o_data_a = 16'b1110110000010000;
            14'h2d26: o_data_a = 16'b0000000000001110;
            14'h2d27: o_data_a = 16'b1110001100001000;
            14'h2d28: o_data_a = 16'b0010110100101100;
            14'h2d29: o_data_a = 16'b1110110000010000;
            14'h2d2a: o_data_a = 16'b0000000001011111;
            14'h2d2b: o_data_a = 16'b1110101010000111;
            14'h2d2c: o_data_a = 16'b0000000000000000;
            14'h2d2d: o_data_a = 16'b1111110010101000;
            14'h2d2e: o_data_a = 16'b1111110000010000;
            14'h2d2f: o_data_a = 16'b0000000000000101;
            14'h2d30: o_data_a = 16'b1110001100001000;
            14'h2d31: o_data_a = 16'b0000000000110011;
            14'h2d32: o_data_a = 16'b1110110000010000;
            14'h2d33: o_data_a = 16'b0000000000000000;
            14'h2d34: o_data_a = 16'b1111110111101000;
            14'h2d35: o_data_a = 16'b1110110010100000;
            14'h2d36: o_data_a = 16'b1110001100001000;
            14'h2d37: o_data_a = 16'b0000000000011110;
            14'h2d38: o_data_a = 16'b1110110000010000;
            14'h2d39: o_data_a = 16'b0000000000000000;
            14'h2d3a: o_data_a = 16'b1111110111101000;
            14'h2d3b: o_data_a = 16'b1110110010100000;
            14'h2d3c: o_data_a = 16'b1110001100001000;
            14'h2d3d: o_data_a = 16'b0000000000110011;
            14'h2d3e: o_data_a = 16'b1110110000010000;
            14'h2d3f: o_data_a = 16'b0000000000000000;
            14'h2d40: o_data_a = 16'b1111110111101000;
            14'h2d41: o_data_a = 16'b1110110010100000;
            14'h2d42: o_data_a = 16'b1110001100001000;
            14'h2d43: o_data_a = 16'b0000000000110000;
            14'h2d44: o_data_a = 16'b1110110000010000;
            14'h2d45: o_data_a = 16'b0000000000000000;
            14'h2d46: o_data_a = 16'b1111110111101000;
            14'h2d47: o_data_a = 16'b1110110010100000;
            14'h2d48: o_data_a = 16'b1110001100001000;
            14'h2d49: o_data_a = 16'b0000000000110000;
            14'h2d4a: o_data_a = 16'b1110110000010000;
            14'h2d4b: o_data_a = 16'b0000000000000000;
            14'h2d4c: o_data_a = 16'b1111110111101000;
            14'h2d4d: o_data_a = 16'b1110110010100000;
            14'h2d4e: o_data_a = 16'b1110001100001000;
            14'h2d4f: o_data_a = 16'b0000000000011100;
            14'h2d50: o_data_a = 16'b1110110000010000;
            14'h2d51: o_data_a = 16'b0000000000000000;
            14'h2d52: o_data_a = 16'b1111110111101000;
            14'h2d53: o_data_a = 16'b1110110010100000;
            14'h2d54: o_data_a = 16'b1110001100001000;
            14'h2d55: o_data_a = 16'b0000000000110000;
            14'h2d56: o_data_a = 16'b1110110000010000;
            14'h2d57: o_data_a = 16'b0000000000000000;
            14'h2d58: o_data_a = 16'b1111110111101000;
            14'h2d59: o_data_a = 16'b1110110010100000;
            14'h2d5a: o_data_a = 16'b1110001100001000;
            14'h2d5b: o_data_a = 16'b0000000000110000;
            14'h2d5c: o_data_a = 16'b1110110000010000;
            14'h2d5d: o_data_a = 16'b0000000000000000;
            14'h2d5e: o_data_a = 16'b1111110111101000;
            14'h2d5f: o_data_a = 16'b1110110010100000;
            14'h2d60: o_data_a = 16'b1110001100001000;
            14'h2d61: o_data_a = 16'b0000000000110011;
            14'h2d62: o_data_a = 16'b1110110000010000;
            14'h2d63: o_data_a = 16'b0000000000000000;
            14'h2d64: o_data_a = 16'b1111110111101000;
            14'h2d65: o_data_a = 16'b1110110010100000;
            14'h2d66: o_data_a = 16'b1110001100001000;
            14'h2d67: o_data_a = 16'b0000000000011110;
            14'h2d68: o_data_a = 16'b1110110000010000;
            14'h2d69: o_data_a = 16'b0000000000000000;
            14'h2d6a: o_data_a = 16'b1111110111101000;
            14'h2d6b: o_data_a = 16'b1110110010100000;
            14'h2d6c: o_data_a = 16'b1110001100001000;
            14'h2d6d: o_data_a = 16'b0000000000000000;
            14'h2d6e: o_data_a = 16'b1111110111001000;
            14'h2d6f: o_data_a = 16'b1111110010100000;
            14'h2d70: o_data_a = 16'b1110101010001000;
            14'h2d71: o_data_a = 16'b0000000000000000;
            14'h2d72: o_data_a = 16'b1111110111001000;
            14'h2d73: o_data_a = 16'b1111110010100000;
            14'h2d74: o_data_a = 16'b1110101010001000;
            14'h2d75: o_data_a = 16'b0000000000001100;
            14'h2d76: o_data_a = 16'b1110110000010000;
            14'h2d77: o_data_a = 16'b0000000000001101;
            14'h2d78: o_data_a = 16'b1110001100001000;
            14'h2d79: o_data_a = 16'b0100010110110011;
            14'h2d7a: o_data_a = 16'b1110110000010000;
            14'h2d7b: o_data_a = 16'b0000000000001110;
            14'h2d7c: o_data_a = 16'b1110001100001000;
            14'h2d7d: o_data_a = 16'b0010110110000001;
            14'h2d7e: o_data_a = 16'b1110110000010000;
            14'h2d7f: o_data_a = 16'b0000000001011111;
            14'h2d80: o_data_a = 16'b1110101010000111;
            14'h2d81: o_data_a = 16'b0000000000000000;
            14'h2d82: o_data_a = 16'b1111110010101000;
            14'h2d83: o_data_a = 16'b1111110000010000;
            14'h2d84: o_data_a = 16'b0000000000000101;
            14'h2d85: o_data_a = 16'b1110001100001000;
            14'h2d86: o_data_a = 16'b0000000000110100;
            14'h2d87: o_data_a = 16'b1110110000010000;
            14'h2d88: o_data_a = 16'b0000000000000000;
            14'h2d89: o_data_a = 16'b1111110111101000;
            14'h2d8a: o_data_a = 16'b1110110010100000;
            14'h2d8b: o_data_a = 16'b1110001100001000;
            14'h2d8c: o_data_a = 16'b0000000000010000;
            14'h2d8d: o_data_a = 16'b1110110000010000;
            14'h2d8e: o_data_a = 16'b0000000000000000;
            14'h2d8f: o_data_a = 16'b1111110111101000;
            14'h2d90: o_data_a = 16'b1110110010100000;
            14'h2d91: o_data_a = 16'b1110001100001000;
            14'h2d92: o_data_a = 16'b0000000000011000;
            14'h2d93: o_data_a = 16'b1110110000010000;
            14'h2d94: o_data_a = 16'b0000000000000000;
            14'h2d95: o_data_a = 16'b1111110111101000;
            14'h2d96: o_data_a = 16'b1110110010100000;
            14'h2d97: o_data_a = 16'b1110001100001000;
            14'h2d98: o_data_a = 16'b0000000000011100;
            14'h2d99: o_data_a = 16'b1110110000010000;
            14'h2d9a: o_data_a = 16'b0000000000000000;
            14'h2d9b: o_data_a = 16'b1111110111101000;
            14'h2d9c: o_data_a = 16'b1110110010100000;
            14'h2d9d: o_data_a = 16'b1110001100001000;
            14'h2d9e: o_data_a = 16'b0000000000011010;
            14'h2d9f: o_data_a = 16'b1110110000010000;
            14'h2da0: o_data_a = 16'b0000000000000000;
            14'h2da1: o_data_a = 16'b1111110111101000;
            14'h2da2: o_data_a = 16'b1110110010100000;
            14'h2da3: o_data_a = 16'b1110001100001000;
            14'h2da4: o_data_a = 16'b0000000000011001;
            14'h2da5: o_data_a = 16'b1110110000010000;
            14'h2da6: o_data_a = 16'b0000000000000000;
            14'h2da7: o_data_a = 16'b1111110111101000;
            14'h2da8: o_data_a = 16'b1110110010100000;
            14'h2da9: o_data_a = 16'b1110001100001000;
            14'h2daa: o_data_a = 16'b0000000000111111;
            14'h2dab: o_data_a = 16'b1110110000010000;
            14'h2dac: o_data_a = 16'b0000000000000000;
            14'h2dad: o_data_a = 16'b1111110111101000;
            14'h2dae: o_data_a = 16'b1110110010100000;
            14'h2daf: o_data_a = 16'b1110001100001000;
            14'h2db0: o_data_a = 16'b0000000000011000;
            14'h2db1: o_data_a = 16'b1110110000010000;
            14'h2db2: o_data_a = 16'b0000000000000000;
            14'h2db3: o_data_a = 16'b1111110111101000;
            14'h2db4: o_data_a = 16'b1110110010100000;
            14'h2db5: o_data_a = 16'b1110001100001000;
            14'h2db6: o_data_a = 16'b0000000000011000;
            14'h2db7: o_data_a = 16'b1110110000010000;
            14'h2db8: o_data_a = 16'b0000000000000000;
            14'h2db9: o_data_a = 16'b1111110111101000;
            14'h2dba: o_data_a = 16'b1110110010100000;
            14'h2dbb: o_data_a = 16'b1110001100001000;
            14'h2dbc: o_data_a = 16'b0000000000111100;
            14'h2dbd: o_data_a = 16'b1110110000010000;
            14'h2dbe: o_data_a = 16'b0000000000000000;
            14'h2dbf: o_data_a = 16'b1111110111101000;
            14'h2dc0: o_data_a = 16'b1110110010100000;
            14'h2dc1: o_data_a = 16'b1110001100001000;
            14'h2dc2: o_data_a = 16'b0000000000000000;
            14'h2dc3: o_data_a = 16'b1111110111001000;
            14'h2dc4: o_data_a = 16'b1111110010100000;
            14'h2dc5: o_data_a = 16'b1110101010001000;
            14'h2dc6: o_data_a = 16'b0000000000000000;
            14'h2dc7: o_data_a = 16'b1111110111001000;
            14'h2dc8: o_data_a = 16'b1111110010100000;
            14'h2dc9: o_data_a = 16'b1110101010001000;
            14'h2dca: o_data_a = 16'b0000000000001100;
            14'h2dcb: o_data_a = 16'b1110110000010000;
            14'h2dcc: o_data_a = 16'b0000000000001101;
            14'h2dcd: o_data_a = 16'b1110001100001000;
            14'h2dce: o_data_a = 16'b0100010110110011;
            14'h2dcf: o_data_a = 16'b1110110000010000;
            14'h2dd0: o_data_a = 16'b0000000000001110;
            14'h2dd1: o_data_a = 16'b1110001100001000;
            14'h2dd2: o_data_a = 16'b0010110111010110;
            14'h2dd3: o_data_a = 16'b1110110000010000;
            14'h2dd4: o_data_a = 16'b0000000001011111;
            14'h2dd5: o_data_a = 16'b1110101010000111;
            14'h2dd6: o_data_a = 16'b0000000000000000;
            14'h2dd7: o_data_a = 16'b1111110010101000;
            14'h2dd8: o_data_a = 16'b1111110000010000;
            14'h2dd9: o_data_a = 16'b0000000000000101;
            14'h2dda: o_data_a = 16'b1110001100001000;
            14'h2ddb: o_data_a = 16'b0000000000110101;
            14'h2ddc: o_data_a = 16'b1110110000010000;
            14'h2ddd: o_data_a = 16'b0000000000000000;
            14'h2dde: o_data_a = 16'b1111110111101000;
            14'h2ddf: o_data_a = 16'b1110110010100000;
            14'h2de0: o_data_a = 16'b1110001100001000;
            14'h2de1: o_data_a = 16'b0000000000111111;
            14'h2de2: o_data_a = 16'b1110110000010000;
            14'h2de3: o_data_a = 16'b0000000000000000;
            14'h2de4: o_data_a = 16'b1111110111101000;
            14'h2de5: o_data_a = 16'b1110110010100000;
            14'h2de6: o_data_a = 16'b1110001100001000;
            14'h2de7: o_data_a = 16'b0000000000000011;
            14'h2de8: o_data_a = 16'b1110110000010000;
            14'h2de9: o_data_a = 16'b0000000000000000;
            14'h2dea: o_data_a = 16'b1111110111101000;
            14'h2deb: o_data_a = 16'b1110110010100000;
            14'h2dec: o_data_a = 16'b1110001100001000;
            14'h2ded: o_data_a = 16'b0000000000000011;
            14'h2dee: o_data_a = 16'b1110110000010000;
            14'h2def: o_data_a = 16'b0000000000000000;
            14'h2df0: o_data_a = 16'b1111110111101000;
            14'h2df1: o_data_a = 16'b1110110010100000;
            14'h2df2: o_data_a = 16'b1110001100001000;
            14'h2df3: o_data_a = 16'b0000000000011111;
            14'h2df4: o_data_a = 16'b1110110000010000;
            14'h2df5: o_data_a = 16'b0000000000000000;
            14'h2df6: o_data_a = 16'b1111110111101000;
            14'h2df7: o_data_a = 16'b1110110010100000;
            14'h2df8: o_data_a = 16'b1110001100001000;
            14'h2df9: o_data_a = 16'b0000000000110000;
            14'h2dfa: o_data_a = 16'b1110110000010000;
            14'h2dfb: o_data_a = 16'b0000000000000000;
            14'h2dfc: o_data_a = 16'b1111110111101000;
            14'h2dfd: o_data_a = 16'b1110110010100000;
            14'h2dfe: o_data_a = 16'b1110001100001000;
            14'h2dff: o_data_a = 16'b0000000000110000;
            14'h2e00: o_data_a = 16'b1110110000010000;
            14'h2e01: o_data_a = 16'b0000000000000000;
            14'h2e02: o_data_a = 16'b1111110111101000;
            14'h2e03: o_data_a = 16'b1110110010100000;
            14'h2e04: o_data_a = 16'b1110001100001000;
            14'h2e05: o_data_a = 16'b0000000000110000;
            14'h2e06: o_data_a = 16'b1110110000010000;
            14'h2e07: o_data_a = 16'b0000000000000000;
            14'h2e08: o_data_a = 16'b1111110111101000;
            14'h2e09: o_data_a = 16'b1110110010100000;
            14'h2e0a: o_data_a = 16'b1110001100001000;
            14'h2e0b: o_data_a = 16'b0000000000110011;
            14'h2e0c: o_data_a = 16'b1110110000010000;
            14'h2e0d: o_data_a = 16'b0000000000000000;
            14'h2e0e: o_data_a = 16'b1111110111101000;
            14'h2e0f: o_data_a = 16'b1110110010100000;
            14'h2e10: o_data_a = 16'b1110001100001000;
            14'h2e11: o_data_a = 16'b0000000000011110;
            14'h2e12: o_data_a = 16'b1110110000010000;
            14'h2e13: o_data_a = 16'b0000000000000000;
            14'h2e14: o_data_a = 16'b1111110111101000;
            14'h2e15: o_data_a = 16'b1110110010100000;
            14'h2e16: o_data_a = 16'b1110001100001000;
            14'h2e17: o_data_a = 16'b0000000000000000;
            14'h2e18: o_data_a = 16'b1111110111001000;
            14'h2e19: o_data_a = 16'b1111110010100000;
            14'h2e1a: o_data_a = 16'b1110101010001000;
            14'h2e1b: o_data_a = 16'b0000000000000000;
            14'h2e1c: o_data_a = 16'b1111110111001000;
            14'h2e1d: o_data_a = 16'b1111110010100000;
            14'h2e1e: o_data_a = 16'b1110101010001000;
            14'h2e1f: o_data_a = 16'b0000000000001100;
            14'h2e20: o_data_a = 16'b1110110000010000;
            14'h2e21: o_data_a = 16'b0000000000001101;
            14'h2e22: o_data_a = 16'b1110001100001000;
            14'h2e23: o_data_a = 16'b0100010110110011;
            14'h2e24: o_data_a = 16'b1110110000010000;
            14'h2e25: o_data_a = 16'b0000000000001110;
            14'h2e26: o_data_a = 16'b1110001100001000;
            14'h2e27: o_data_a = 16'b0010111000101011;
            14'h2e28: o_data_a = 16'b1110110000010000;
            14'h2e29: o_data_a = 16'b0000000001011111;
            14'h2e2a: o_data_a = 16'b1110101010000111;
            14'h2e2b: o_data_a = 16'b0000000000000000;
            14'h2e2c: o_data_a = 16'b1111110010101000;
            14'h2e2d: o_data_a = 16'b1111110000010000;
            14'h2e2e: o_data_a = 16'b0000000000000101;
            14'h2e2f: o_data_a = 16'b1110001100001000;
            14'h2e30: o_data_a = 16'b0000000000110110;
            14'h2e31: o_data_a = 16'b1110110000010000;
            14'h2e32: o_data_a = 16'b0000000000000000;
            14'h2e33: o_data_a = 16'b1111110111101000;
            14'h2e34: o_data_a = 16'b1110110010100000;
            14'h2e35: o_data_a = 16'b1110001100001000;
            14'h2e36: o_data_a = 16'b0000000000011100;
            14'h2e37: o_data_a = 16'b1110110000010000;
            14'h2e38: o_data_a = 16'b0000000000000000;
            14'h2e39: o_data_a = 16'b1111110111101000;
            14'h2e3a: o_data_a = 16'b1110110010100000;
            14'h2e3b: o_data_a = 16'b1110001100001000;
            14'h2e3c: o_data_a = 16'b0000000000000110;
            14'h2e3d: o_data_a = 16'b1110110000010000;
            14'h2e3e: o_data_a = 16'b0000000000000000;
            14'h2e3f: o_data_a = 16'b1111110111101000;
            14'h2e40: o_data_a = 16'b1110110010100000;
            14'h2e41: o_data_a = 16'b1110001100001000;
            14'h2e42: o_data_a = 16'b0000000000000011;
            14'h2e43: o_data_a = 16'b1110110000010000;
            14'h2e44: o_data_a = 16'b0000000000000000;
            14'h2e45: o_data_a = 16'b1111110111101000;
            14'h2e46: o_data_a = 16'b1110110010100000;
            14'h2e47: o_data_a = 16'b1110001100001000;
            14'h2e48: o_data_a = 16'b0000000000000011;
            14'h2e49: o_data_a = 16'b1110110000010000;
            14'h2e4a: o_data_a = 16'b0000000000000000;
            14'h2e4b: o_data_a = 16'b1111110111101000;
            14'h2e4c: o_data_a = 16'b1110110010100000;
            14'h2e4d: o_data_a = 16'b1110001100001000;
            14'h2e4e: o_data_a = 16'b0000000000011111;
            14'h2e4f: o_data_a = 16'b1110110000010000;
            14'h2e50: o_data_a = 16'b0000000000000000;
            14'h2e51: o_data_a = 16'b1111110111101000;
            14'h2e52: o_data_a = 16'b1110110010100000;
            14'h2e53: o_data_a = 16'b1110001100001000;
            14'h2e54: o_data_a = 16'b0000000000110011;
            14'h2e55: o_data_a = 16'b1110110000010000;
            14'h2e56: o_data_a = 16'b0000000000000000;
            14'h2e57: o_data_a = 16'b1111110111101000;
            14'h2e58: o_data_a = 16'b1110110010100000;
            14'h2e59: o_data_a = 16'b1110001100001000;
            14'h2e5a: o_data_a = 16'b0000000000110011;
            14'h2e5b: o_data_a = 16'b1110110000010000;
            14'h2e5c: o_data_a = 16'b0000000000000000;
            14'h2e5d: o_data_a = 16'b1111110111101000;
            14'h2e5e: o_data_a = 16'b1110110010100000;
            14'h2e5f: o_data_a = 16'b1110001100001000;
            14'h2e60: o_data_a = 16'b0000000000110011;
            14'h2e61: o_data_a = 16'b1110110000010000;
            14'h2e62: o_data_a = 16'b0000000000000000;
            14'h2e63: o_data_a = 16'b1111110111101000;
            14'h2e64: o_data_a = 16'b1110110010100000;
            14'h2e65: o_data_a = 16'b1110001100001000;
            14'h2e66: o_data_a = 16'b0000000000011110;
            14'h2e67: o_data_a = 16'b1110110000010000;
            14'h2e68: o_data_a = 16'b0000000000000000;
            14'h2e69: o_data_a = 16'b1111110111101000;
            14'h2e6a: o_data_a = 16'b1110110010100000;
            14'h2e6b: o_data_a = 16'b1110001100001000;
            14'h2e6c: o_data_a = 16'b0000000000000000;
            14'h2e6d: o_data_a = 16'b1111110111001000;
            14'h2e6e: o_data_a = 16'b1111110010100000;
            14'h2e6f: o_data_a = 16'b1110101010001000;
            14'h2e70: o_data_a = 16'b0000000000000000;
            14'h2e71: o_data_a = 16'b1111110111001000;
            14'h2e72: o_data_a = 16'b1111110010100000;
            14'h2e73: o_data_a = 16'b1110101010001000;
            14'h2e74: o_data_a = 16'b0000000000001100;
            14'h2e75: o_data_a = 16'b1110110000010000;
            14'h2e76: o_data_a = 16'b0000000000001101;
            14'h2e77: o_data_a = 16'b1110001100001000;
            14'h2e78: o_data_a = 16'b0100010110110011;
            14'h2e79: o_data_a = 16'b1110110000010000;
            14'h2e7a: o_data_a = 16'b0000000000001110;
            14'h2e7b: o_data_a = 16'b1110001100001000;
            14'h2e7c: o_data_a = 16'b0010111010000000;
            14'h2e7d: o_data_a = 16'b1110110000010000;
            14'h2e7e: o_data_a = 16'b0000000001011111;
            14'h2e7f: o_data_a = 16'b1110101010000111;
            14'h2e80: o_data_a = 16'b0000000000000000;
            14'h2e81: o_data_a = 16'b1111110010101000;
            14'h2e82: o_data_a = 16'b1111110000010000;
            14'h2e83: o_data_a = 16'b0000000000000101;
            14'h2e84: o_data_a = 16'b1110001100001000;
            14'h2e85: o_data_a = 16'b0000000000110111;
            14'h2e86: o_data_a = 16'b1110110000010000;
            14'h2e87: o_data_a = 16'b0000000000000000;
            14'h2e88: o_data_a = 16'b1111110111101000;
            14'h2e89: o_data_a = 16'b1110110010100000;
            14'h2e8a: o_data_a = 16'b1110001100001000;
            14'h2e8b: o_data_a = 16'b0000000000111111;
            14'h2e8c: o_data_a = 16'b1110110000010000;
            14'h2e8d: o_data_a = 16'b0000000000000000;
            14'h2e8e: o_data_a = 16'b1111110111101000;
            14'h2e8f: o_data_a = 16'b1110110010100000;
            14'h2e90: o_data_a = 16'b1110001100001000;
            14'h2e91: o_data_a = 16'b0000000000110001;
            14'h2e92: o_data_a = 16'b1110110000010000;
            14'h2e93: o_data_a = 16'b0000000000000000;
            14'h2e94: o_data_a = 16'b1111110111101000;
            14'h2e95: o_data_a = 16'b1110110010100000;
            14'h2e96: o_data_a = 16'b1110001100001000;
            14'h2e97: o_data_a = 16'b0000000000110000;
            14'h2e98: o_data_a = 16'b1110110000010000;
            14'h2e99: o_data_a = 16'b0000000000000000;
            14'h2e9a: o_data_a = 16'b1111110111101000;
            14'h2e9b: o_data_a = 16'b1110110010100000;
            14'h2e9c: o_data_a = 16'b1110001100001000;
            14'h2e9d: o_data_a = 16'b0000000000110000;
            14'h2e9e: o_data_a = 16'b1110110000010000;
            14'h2e9f: o_data_a = 16'b0000000000000000;
            14'h2ea0: o_data_a = 16'b1111110111101000;
            14'h2ea1: o_data_a = 16'b1110110010100000;
            14'h2ea2: o_data_a = 16'b1110001100001000;
            14'h2ea3: o_data_a = 16'b0000000000011000;
            14'h2ea4: o_data_a = 16'b1110110000010000;
            14'h2ea5: o_data_a = 16'b0000000000000000;
            14'h2ea6: o_data_a = 16'b1111110111101000;
            14'h2ea7: o_data_a = 16'b1110110010100000;
            14'h2ea8: o_data_a = 16'b1110001100001000;
            14'h2ea9: o_data_a = 16'b0000000000001100;
            14'h2eaa: o_data_a = 16'b1110110000010000;
            14'h2eab: o_data_a = 16'b0000000000000000;
            14'h2eac: o_data_a = 16'b1111110111101000;
            14'h2ead: o_data_a = 16'b1110110010100000;
            14'h2eae: o_data_a = 16'b1110001100001000;
            14'h2eaf: o_data_a = 16'b0000000000001100;
            14'h2eb0: o_data_a = 16'b1110110000010000;
            14'h2eb1: o_data_a = 16'b0000000000000000;
            14'h2eb2: o_data_a = 16'b1111110111101000;
            14'h2eb3: o_data_a = 16'b1110110010100000;
            14'h2eb4: o_data_a = 16'b1110001100001000;
            14'h2eb5: o_data_a = 16'b0000000000001100;
            14'h2eb6: o_data_a = 16'b1110110000010000;
            14'h2eb7: o_data_a = 16'b0000000000000000;
            14'h2eb8: o_data_a = 16'b1111110111101000;
            14'h2eb9: o_data_a = 16'b1110110010100000;
            14'h2eba: o_data_a = 16'b1110001100001000;
            14'h2ebb: o_data_a = 16'b0000000000001100;
            14'h2ebc: o_data_a = 16'b1110110000010000;
            14'h2ebd: o_data_a = 16'b0000000000000000;
            14'h2ebe: o_data_a = 16'b1111110111101000;
            14'h2ebf: o_data_a = 16'b1110110010100000;
            14'h2ec0: o_data_a = 16'b1110001100001000;
            14'h2ec1: o_data_a = 16'b0000000000000000;
            14'h2ec2: o_data_a = 16'b1111110111001000;
            14'h2ec3: o_data_a = 16'b1111110010100000;
            14'h2ec4: o_data_a = 16'b1110101010001000;
            14'h2ec5: o_data_a = 16'b0000000000000000;
            14'h2ec6: o_data_a = 16'b1111110111001000;
            14'h2ec7: o_data_a = 16'b1111110010100000;
            14'h2ec8: o_data_a = 16'b1110101010001000;
            14'h2ec9: o_data_a = 16'b0000000000001100;
            14'h2eca: o_data_a = 16'b1110110000010000;
            14'h2ecb: o_data_a = 16'b0000000000001101;
            14'h2ecc: o_data_a = 16'b1110001100001000;
            14'h2ecd: o_data_a = 16'b0100010110110011;
            14'h2ece: o_data_a = 16'b1110110000010000;
            14'h2ecf: o_data_a = 16'b0000000000001110;
            14'h2ed0: o_data_a = 16'b1110001100001000;
            14'h2ed1: o_data_a = 16'b0010111011010101;
            14'h2ed2: o_data_a = 16'b1110110000010000;
            14'h2ed3: o_data_a = 16'b0000000001011111;
            14'h2ed4: o_data_a = 16'b1110101010000111;
            14'h2ed5: o_data_a = 16'b0000000000000000;
            14'h2ed6: o_data_a = 16'b1111110010101000;
            14'h2ed7: o_data_a = 16'b1111110000010000;
            14'h2ed8: o_data_a = 16'b0000000000000101;
            14'h2ed9: o_data_a = 16'b1110001100001000;
            14'h2eda: o_data_a = 16'b0000000000111000;
            14'h2edb: o_data_a = 16'b1110110000010000;
            14'h2edc: o_data_a = 16'b0000000000000000;
            14'h2edd: o_data_a = 16'b1111110111101000;
            14'h2ede: o_data_a = 16'b1110110010100000;
            14'h2edf: o_data_a = 16'b1110001100001000;
            14'h2ee0: o_data_a = 16'b0000000000011110;
            14'h2ee1: o_data_a = 16'b1110110000010000;
            14'h2ee2: o_data_a = 16'b0000000000000000;
            14'h2ee3: o_data_a = 16'b1111110111101000;
            14'h2ee4: o_data_a = 16'b1110110010100000;
            14'h2ee5: o_data_a = 16'b1110001100001000;
            14'h2ee6: o_data_a = 16'b0000000000110011;
            14'h2ee7: o_data_a = 16'b1110110000010000;
            14'h2ee8: o_data_a = 16'b0000000000000000;
            14'h2ee9: o_data_a = 16'b1111110111101000;
            14'h2eea: o_data_a = 16'b1110110010100000;
            14'h2eeb: o_data_a = 16'b1110001100001000;
            14'h2eec: o_data_a = 16'b0000000000110011;
            14'h2eed: o_data_a = 16'b1110110000010000;
            14'h2eee: o_data_a = 16'b0000000000000000;
            14'h2eef: o_data_a = 16'b1111110111101000;
            14'h2ef0: o_data_a = 16'b1110110010100000;
            14'h2ef1: o_data_a = 16'b1110001100001000;
            14'h2ef2: o_data_a = 16'b0000000000110011;
            14'h2ef3: o_data_a = 16'b1110110000010000;
            14'h2ef4: o_data_a = 16'b0000000000000000;
            14'h2ef5: o_data_a = 16'b1111110111101000;
            14'h2ef6: o_data_a = 16'b1110110010100000;
            14'h2ef7: o_data_a = 16'b1110001100001000;
            14'h2ef8: o_data_a = 16'b0000000000011110;
            14'h2ef9: o_data_a = 16'b1110110000010000;
            14'h2efa: o_data_a = 16'b0000000000000000;
            14'h2efb: o_data_a = 16'b1111110111101000;
            14'h2efc: o_data_a = 16'b1110110010100000;
            14'h2efd: o_data_a = 16'b1110001100001000;
            14'h2efe: o_data_a = 16'b0000000000110011;
            14'h2eff: o_data_a = 16'b1110110000010000;
            14'h2f00: o_data_a = 16'b0000000000000000;
            14'h2f01: o_data_a = 16'b1111110111101000;
            14'h2f02: o_data_a = 16'b1110110010100000;
            14'h2f03: o_data_a = 16'b1110001100001000;
            14'h2f04: o_data_a = 16'b0000000000110011;
            14'h2f05: o_data_a = 16'b1110110000010000;
            14'h2f06: o_data_a = 16'b0000000000000000;
            14'h2f07: o_data_a = 16'b1111110111101000;
            14'h2f08: o_data_a = 16'b1110110010100000;
            14'h2f09: o_data_a = 16'b1110001100001000;
            14'h2f0a: o_data_a = 16'b0000000000110011;
            14'h2f0b: o_data_a = 16'b1110110000010000;
            14'h2f0c: o_data_a = 16'b0000000000000000;
            14'h2f0d: o_data_a = 16'b1111110111101000;
            14'h2f0e: o_data_a = 16'b1110110010100000;
            14'h2f0f: o_data_a = 16'b1110001100001000;
            14'h2f10: o_data_a = 16'b0000000000011110;
            14'h2f11: o_data_a = 16'b1110110000010000;
            14'h2f12: o_data_a = 16'b0000000000000000;
            14'h2f13: o_data_a = 16'b1111110111101000;
            14'h2f14: o_data_a = 16'b1110110010100000;
            14'h2f15: o_data_a = 16'b1110001100001000;
            14'h2f16: o_data_a = 16'b0000000000000000;
            14'h2f17: o_data_a = 16'b1111110111001000;
            14'h2f18: o_data_a = 16'b1111110010100000;
            14'h2f19: o_data_a = 16'b1110101010001000;
            14'h2f1a: o_data_a = 16'b0000000000000000;
            14'h2f1b: o_data_a = 16'b1111110111001000;
            14'h2f1c: o_data_a = 16'b1111110010100000;
            14'h2f1d: o_data_a = 16'b1110101010001000;
            14'h2f1e: o_data_a = 16'b0000000000001100;
            14'h2f1f: o_data_a = 16'b1110110000010000;
            14'h2f20: o_data_a = 16'b0000000000001101;
            14'h2f21: o_data_a = 16'b1110001100001000;
            14'h2f22: o_data_a = 16'b0100010110110011;
            14'h2f23: o_data_a = 16'b1110110000010000;
            14'h2f24: o_data_a = 16'b0000000000001110;
            14'h2f25: o_data_a = 16'b1110001100001000;
            14'h2f26: o_data_a = 16'b0010111100101010;
            14'h2f27: o_data_a = 16'b1110110000010000;
            14'h2f28: o_data_a = 16'b0000000001011111;
            14'h2f29: o_data_a = 16'b1110101010000111;
            14'h2f2a: o_data_a = 16'b0000000000000000;
            14'h2f2b: o_data_a = 16'b1111110010101000;
            14'h2f2c: o_data_a = 16'b1111110000010000;
            14'h2f2d: o_data_a = 16'b0000000000000101;
            14'h2f2e: o_data_a = 16'b1110001100001000;
            14'h2f2f: o_data_a = 16'b0000000000111001;
            14'h2f30: o_data_a = 16'b1110110000010000;
            14'h2f31: o_data_a = 16'b0000000000000000;
            14'h2f32: o_data_a = 16'b1111110111101000;
            14'h2f33: o_data_a = 16'b1110110010100000;
            14'h2f34: o_data_a = 16'b1110001100001000;
            14'h2f35: o_data_a = 16'b0000000000011110;
            14'h2f36: o_data_a = 16'b1110110000010000;
            14'h2f37: o_data_a = 16'b0000000000000000;
            14'h2f38: o_data_a = 16'b1111110111101000;
            14'h2f39: o_data_a = 16'b1110110010100000;
            14'h2f3a: o_data_a = 16'b1110001100001000;
            14'h2f3b: o_data_a = 16'b0000000000110011;
            14'h2f3c: o_data_a = 16'b1110110000010000;
            14'h2f3d: o_data_a = 16'b0000000000000000;
            14'h2f3e: o_data_a = 16'b1111110111101000;
            14'h2f3f: o_data_a = 16'b1110110010100000;
            14'h2f40: o_data_a = 16'b1110001100001000;
            14'h2f41: o_data_a = 16'b0000000000110011;
            14'h2f42: o_data_a = 16'b1110110000010000;
            14'h2f43: o_data_a = 16'b0000000000000000;
            14'h2f44: o_data_a = 16'b1111110111101000;
            14'h2f45: o_data_a = 16'b1110110010100000;
            14'h2f46: o_data_a = 16'b1110001100001000;
            14'h2f47: o_data_a = 16'b0000000000110011;
            14'h2f48: o_data_a = 16'b1110110000010000;
            14'h2f49: o_data_a = 16'b0000000000000000;
            14'h2f4a: o_data_a = 16'b1111110111101000;
            14'h2f4b: o_data_a = 16'b1110110010100000;
            14'h2f4c: o_data_a = 16'b1110001100001000;
            14'h2f4d: o_data_a = 16'b0000000000111110;
            14'h2f4e: o_data_a = 16'b1110110000010000;
            14'h2f4f: o_data_a = 16'b0000000000000000;
            14'h2f50: o_data_a = 16'b1111110111101000;
            14'h2f51: o_data_a = 16'b1110110010100000;
            14'h2f52: o_data_a = 16'b1110001100001000;
            14'h2f53: o_data_a = 16'b0000000000110000;
            14'h2f54: o_data_a = 16'b1110110000010000;
            14'h2f55: o_data_a = 16'b0000000000000000;
            14'h2f56: o_data_a = 16'b1111110111101000;
            14'h2f57: o_data_a = 16'b1110110010100000;
            14'h2f58: o_data_a = 16'b1110001100001000;
            14'h2f59: o_data_a = 16'b0000000000110000;
            14'h2f5a: o_data_a = 16'b1110110000010000;
            14'h2f5b: o_data_a = 16'b0000000000000000;
            14'h2f5c: o_data_a = 16'b1111110111101000;
            14'h2f5d: o_data_a = 16'b1110110010100000;
            14'h2f5e: o_data_a = 16'b1110001100001000;
            14'h2f5f: o_data_a = 16'b0000000000011000;
            14'h2f60: o_data_a = 16'b1110110000010000;
            14'h2f61: o_data_a = 16'b0000000000000000;
            14'h2f62: o_data_a = 16'b1111110111101000;
            14'h2f63: o_data_a = 16'b1110110010100000;
            14'h2f64: o_data_a = 16'b1110001100001000;
            14'h2f65: o_data_a = 16'b0000000000001110;
            14'h2f66: o_data_a = 16'b1110110000010000;
            14'h2f67: o_data_a = 16'b0000000000000000;
            14'h2f68: o_data_a = 16'b1111110111101000;
            14'h2f69: o_data_a = 16'b1110110010100000;
            14'h2f6a: o_data_a = 16'b1110001100001000;
            14'h2f6b: o_data_a = 16'b0000000000000000;
            14'h2f6c: o_data_a = 16'b1111110111001000;
            14'h2f6d: o_data_a = 16'b1111110010100000;
            14'h2f6e: o_data_a = 16'b1110101010001000;
            14'h2f6f: o_data_a = 16'b0000000000000000;
            14'h2f70: o_data_a = 16'b1111110111001000;
            14'h2f71: o_data_a = 16'b1111110010100000;
            14'h2f72: o_data_a = 16'b1110101010001000;
            14'h2f73: o_data_a = 16'b0000000000001100;
            14'h2f74: o_data_a = 16'b1110110000010000;
            14'h2f75: o_data_a = 16'b0000000000001101;
            14'h2f76: o_data_a = 16'b1110001100001000;
            14'h2f77: o_data_a = 16'b0100010110110011;
            14'h2f78: o_data_a = 16'b1110110000010000;
            14'h2f79: o_data_a = 16'b0000000000001110;
            14'h2f7a: o_data_a = 16'b1110001100001000;
            14'h2f7b: o_data_a = 16'b0010111101111111;
            14'h2f7c: o_data_a = 16'b1110110000010000;
            14'h2f7d: o_data_a = 16'b0000000001011111;
            14'h2f7e: o_data_a = 16'b1110101010000111;
            14'h2f7f: o_data_a = 16'b0000000000000000;
            14'h2f80: o_data_a = 16'b1111110010101000;
            14'h2f81: o_data_a = 16'b1111110000010000;
            14'h2f82: o_data_a = 16'b0000000000000101;
            14'h2f83: o_data_a = 16'b1110001100001000;
            14'h2f84: o_data_a = 16'b0000000000111010;
            14'h2f85: o_data_a = 16'b1110110000010000;
            14'h2f86: o_data_a = 16'b0000000000000000;
            14'h2f87: o_data_a = 16'b1111110111101000;
            14'h2f88: o_data_a = 16'b1110110010100000;
            14'h2f89: o_data_a = 16'b1110001100001000;
            14'h2f8a: o_data_a = 16'b0000000000000000;
            14'h2f8b: o_data_a = 16'b1111110111001000;
            14'h2f8c: o_data_a = 16'b1111110010100000;
            14'h2f8d: o_data_a = 16'b1110101010001000;
            14'h2f8e: o_data_a = 16'b0000000000000000;
            14'h2f8f: o_data_a = 16'b1111110111001000;
            14'h2f90: o_data_a = 16'b1111110010100000;
            14'h2f91: o_data_a = 16'b1110101010001000;
            14'h2f92: o_data_a = 16'b0000000000001100;
            14'h2f93: o_data_a = 16'b1110110000010000;
            14'h2f94: o_data_a = 16'b0000000000000000;
            14'h2f95: o_data_a = 16'b1111110111101000;
            14'h2f96: o_data_a = 16'b1110110010100000;
            14'h2f97: o_data_a = 16'b1110001100001000;
            14'h2f98: o_data_a = 16'b0000000000001100;
            14'h2f99: o_data_a = 16'b1110110000010000;
            14'h2f9a: o_data_a = 16'b0000000000000000;
            14'h2f9b: o_data_a = 16'b1111110111101000;
            14'h2f9c: o_data_a = 16'b1110110010100000;
            14'h2f9d: o_data_a = 16'b1110001100001000;
            14'h2f9e: o_data_a = 16'b0000000000000000;
            14'h2f9f: o_data_a = 16'b1111110111001000;
            14'h2fa0: o_data_a = 16'b1111110010100000;
            14'h2fa1: o_data_a = 16'b1110101010001000;
            14'h2fa2: o_data_a = 16'b0000000000000000;
            14'h2fa3: o_data_a = 16'b1111110111001000;
            14'h2fa4: o_data_a = 16'b1111110010100000;
            14'h2fa5: o_data_a = 16'b1110101010001000;
            14'h2fa6: o_data_a = 16'b0000000000001100;
            14'h2fa7: o_data_a = 16'b1110110000010000;
            14'h2fa8: o_data_a = 16'b0000000000000000;
            14'h2fa9: o_data_a = 16'b1111110111101000;
            14'h2faa: o_data_a = 16'b1110110010100000;
            14'h2fab: o_data_a = 16'b1110001100001000;
            14'h2fac: o_data_a = 16'b0000000000001100;
            14'h2fad: o_data_a = 16'b1110110000010000;
            14'h2fae: o_data_a = 16'b0000000000000000;
            14'h2faf: o_data_a = 16'b1111110111101000;
            14'h2fb0: o_data_a = 16'b1110110010100000;
            14'h2fb1: o_data_a = 16'b1110001100001000;
            14'h2fb2: o_data_a = 16'b0000000000000000;
            14'h2fb3: o_data_a = 16'b1111110111001000;
            14'h2fb4: o_data_a = 16'b1111110010100000;
            14'h2fb5: o_data_a = 16'b1110101010001000;
            14'h2fb6: o_data_a = 16'b0000000000000000;
            14'h2fb7: o_data_a = 16'b1111110111001000;
            14'h2fb8: o_data_a = 16'b1111110010100000;
            14'h2fb9: o_data_a = 16'b1110101010001000;
            14'h2fba: o_data_a = 16'b0000000000000000;
            14'h2fbb: o_data_a = 16'b1111110111001000;
            14'h2fbc: o_data_a = 16'b1111110010100000;
            14'h2fbd: o_data_a = 16'b1110101010001000;
            14'h2fbe: o_data_a = 16'b0000000000001100;
            14'h2fbf: o_data_a = 16'b1110110000010000;
            14'h2fc0: o_data_a = 16'b0000000000001101;
            14'h2fc1: o_data_a = 16'b1110001100001000;
            14'h2fc2: o_data_a = 16'b0100010110110011;
            14'h2fc3: o_data_a = 16'b1110110000010000;
            14'h2fc4: o_data_a = 16'b0000000000001110;
            14'h2fc5: o_data_a = 16'b1110001100001000;
            14'h2fc6: o_data_a = 16'b0010111111001010;
            14'h2fc7: o_data_a = 16'b1110110000010000;
            14'h2fc8: o_data_a = 16'b0000000001011111;
            14'h2fc9: o_data_a = 16'b1110101010000111;
            14'h2fca: o_data_a = 16'b0000000000000000;
            14'h2fcb: o_data_a = 16'b1111110010101000;
            14'h2fcc: o_data_a = 16'b1111110000010000;
            14'h2fcd: o_data_a = 16'b0000000000000101;
            14'h2fce: o_data_a = 16'b1110001100001000;
            14'h2fcf: o_data_a = 16'b0000000000111011;
            14'h2fd0: o_data_a = 16'b1110110000010000;
            14'h2fd1: o_data_a = 16'b0000000000000000;
            14'h2fd2: o_data_a = 16'b1111110111101000;
            14'h2fd3: o_data_a = 16'b1110110010100000;
            14'h2fd4: o_data_a = 16'b1110001100001000;
            14'h2fd5: o_data_a = 16'b0000000000000000;
            14'h2fd6: o_data_a = 16'b1111110111001000;
            14'h2fd7: o_data_a = 16'b1111110010100000;
            14'h2fd8: o_data_a = 16'b1110101010001000;
            14'h2fd9: o_data_a = 16'b0000000000000000;
            14'h2fda: o_data_a = 16'b1111110111001000;
            14'h2fdb: o_data_a = 16'b1111110010100000;
            14'h2fdc: o_data_a = 16'b1110101010001000;
            14'h2fdd: o_data_a = 16'b0000000000001100;
            14'h2fde: o_data_a = 16'b1110110000010000;
            14'h2fdf: o_data_a = 16'b0000000000000000;
            14'h2fe0: o_data_a = 16'b1111110111101000;
            14'h2fe1: o_data_a = 16'b1110110010100000;
            14'h2fe2: o_data_a = 16'b1110001100001000;
            14'h2fe3: o_data_a = 16'b0000000000001100;
            14'h2fe4: o_data_a = 16'b1110110000010000;
            14'h2fe5: o_data_a = 16'b0000000000000000;
            14'h2fe6: o_data_a = 16'b1111110111101000;
            14'h2fe7: o_data_a = 16'b1110110010100000;
            14'h2fe8: o_data_a = 16'b1110001100001000;
            14'h2fe9: o_data_a = 16'b0000000000000000;
            14'h2fea: o_data_a = 16'b1111110111001000;
            14'h2feb: o_data_a = 16'b1111110010100000;
            14'h2fec: o_data_a = 16'b1110101010001000;
            14'h2fed: o_data_a = 16'b0000000000000000;
            14'h2fee: o_data_a = 16'b1111110111001000;
            14'h2fef: o_data_a = 16'b1111110010100000;
            14'h2ff0: o_data_a = 16'b1110101010001000;
            14'h2ff1: o_data_a = 16'b0000000000001100;
            14'h2ff2: o_data_a = 16'b1110110000010000;
            14'h2ff3: o_data_a = 16'b0000000000000000;
            14'h2ff4: o_data_a = 16'b1111110111101000;
            14'h2ff5: o_data_a = 16'b1110110010100000;
            14'h2ff6: o_data_a = 16'b1110001100001000;
            14'h2ff7: o_data_a = 16'b0000000000001100;
            14'h2ff8: o_data_a = 16'b1110110000010000;
            14'h2ff9: o_data_a = 16'b0000000000000000;
            14'h2ffa: o_data_a = 16'b1111110111101000;
            14'h2ffb: o_data_a = 16'b1110110010100000;
            14'h2ffc: o_data_a = 16'b1110001100001000;
            14'h2ffd: o_data_a = 16'b0000000000000110;
            14'h2ffe: o_data_a = 16'b1110110000010000;
            14'h2fff: o_data_a = 16'b0000000000000000;
            14'h3000: o_data_a = 16'b1111110111101000;
            14'h3001: o_data_a = 16'b1110110010100000;
            14'h3002: o_data_a = 16'b1110001100001000;
            14'h3003: o_data_a = 16'b0000000000000000;
            14'h3004: o_data_a = 16'b1111110111001000;
            14'h3005: o_data_a = 16'b1111110010100000;
            14'h3006: o_data_a = 16'b1110101010001000;
            14'h3007: o_data_a = 16'b0000000000000000;
            14'h3008: o_data_a = 16'b1111110111001000;
            14'h3009: o_data_a = 16'b1111110010100000;
            14'h300a: o_data_a = 16'b1110101010001000;
            14'h300b: o_data_a = 16'b0000000000001100;
            14'h300c: o_data_a = 16'b1110110000010000;
            14'h300d: o_data_a = 16'b0000000000001101;
            14'h300e: o_data_a = 16'b1110001100001000;
            14'h300f: o_data_a = 16'b0100010110110011;
            14'h3010: o_data_a = 16'b1110110000010000;
            14'h3011: o_data_a = 16'b0000000000001110;
            14'h3012: o_data_a = 16'b1110001100001000;
            14'h3013: o_data_a = 16'b0011000000010111;
            14'h3014: o_data_a = 16'b1110110000010000;
            14'h3015: o_data_a = 16'b0000000001011111;
            14'h3016: o_data_a = 16'b1110101010000111;
            14'h3017: o_data_a = 16'b0000000000000000;
            14'h3018: o_data_a = 16'b1111110010101000;
            14'h3019: o_data_a = 16'b1111110000010000;
            14'h301a: o_data_a = 16'b0000000000000101;
            14'h301b: o_data_a = 16'b1110001100001000;
            14'h301c: o_data_a = 16'b0000000000111100;
            14'h301d: o_data_a = 16'b1110110000010000;
            14'h301e: o_data_a = 16'b0000000000000000;
            14'h301f: o_data_a = 16'b1111110111101000;
            14'h3020: o_data_a = 16'b1110110010100000;
            14'h3021: o_data_a = 16'b1110001100001000;
            14'h3022: o_data_a = 16'b0000000000000000;
            14'h3023: o_data_a = 16'b1111110111001000;
            14'h3024: o_data_a = 16'b1111110010100000;
            14'h3025: o_data_a = 16'b1110101010001000;
            14'h3026: o_data_a = 16'b0000000000000000;
            14'h3027: o_data_a = 16'b1111110111001000;
            14'h3028: o_data_a = 16'b1111110010100000;
            14'h3029: o_data_a = 16'b1110101010001000;
            14'h302a: o_data_a = 16'b0000000000011000;
            14'h302b: o_data_a = 16'b1110110000010000;
            14'h302c: o_data_a = 16'b0000000000000000;
            14'h302d: o_data_a = 16'b1111110111101000;
            14'h302e: o_data_a = 16'b1110110010100000;
            14'h302f: o_data_a = 16'b1110001100001000;
            14'h3030: o_data_a = 16'b0000000000001100;
            14'h3031: o_data_a = 16'b1110110000010000;
            14'h3032: o_data_a = 16'b0000000000000000;
            14'h3033: o_data_a = 16'b1111110111101000;
            14'h3034: o_data_a = 16'b1110110010100000;
            14'h3035: o_data_a = 16'b1110001100001000;
            14'h3036: o_data_a = 16'b0000000000000110;
            14'h3037: o_data_a = 16'b1110110000010000;
            14'h3038: o_data_a = 16'b0000000000000000;
            14'h3039: o_data_a = 16'b1111110111101000;
            14'h303a: o_data_a = 16'b1110110010100000;
            14'h303b: o_data_a = 16'b1110001100001000;
            14'h303c: o_data_a = 16'b0000000000000011;
            14'h303d: o_data_a = 16'b1110110000010000;
            14'h303e: o_data_a = 16'b0000000000000000;
            14'h303f: o_data_a = 16'b1111110111101000;
            14'h3040: o_data_a = 16'b1110110010100000;
            14'h3041: o_data_a = 16'b1110001100001000;
            14'h3042: o_data_a = 16'b0000000000000110;
            14'h3043: o_data_a = 16'b1110110000010000;
            14'h3044: o_data_a = 16'b0000000000000000;
            14'h3045: o_data_a = 16'b1111110111101000;
            14'h3046: o_data_a = 16'b1110110010100000;
            14'h3047: o_data_a = 16'b1110001100001000;
            14'h3048: o_data_a = 16'b0000000000001100;
            14'h3049: o_data_a = 16'b1110110000010000;
            14'h304a: o_data_a = 16'b0000000000000000;
            14'h304b: o_data_a = 16'b1111110111101000;
            14'h304c: o_data_a = 16'b1110110010100000;
            14'h304d: o_data_a = 16'b1110001100001000;
            14'h304e: o_data_a = 16'b0000000000011000;
            14'h304f: o_data_a = 16'b1110110000010000;
            14'h3050: o_data_a = 16'b0000000000000000;
            14'h3051: o_data_a = 16'b1111110111101000;
            14'h3052: o_data_a = 16'b1110110010100000;
            14'h3053: o_data_a = 16'b1110001100001000;
            14'h3054: o_data_a = 16'b0000000000000000;
            14'h3055: o_data_a = 16'b1111110111001000;
            14'h3056: o_data_a = 16'b1111110010100000;
            14'h3057: o_data_a = 16'b1110101010001000;
            14'h3058: o_data_a = 16'b0000000000000000;
            14'h3059: o_data_a = 16'b1111110111001000;
            14'h305a: o_data_a = 16'b1111110010100000;
            14'h305b: o_data_a = 16'b1110101010001000;
            14'h305c: o_data_a = 16'b0000000000001100;
            14'h305d: o_data_a = 16'b1110110000010000;
            14'h305e: o_data_a = 16'b0000000000001101;
            14'h305f: o_data_a = 16'b1110001100001000;
            14'h3060: o_data_a = 16'b0100010110110011;
            14'h3061: o_data_a = 16'b1110110000010000;
            14'h3062: o_data_a = 16'b0000000000001110;
            14'h3063: o_data_a = 16'b1110001100001000;
            14'h3064: o_data_a = 16'b0011000001101000;
            14'h3065: o_data_a = 16'b1110110000010000;
            14'h3066: o_data_a = 16'b0000000001011111;
            14'h3067: o_data_a = 16'b1110101010000111;
            14'h3068: o_data_a = 16'b0000000000000000;
            14'h3069: o_data_a = 16'b1111110010101000;
            14'h306a: o_data_a = 16'b1111110000010000;
            14'h306b: o_data_a = 16'b0000000000000101;
            14'h306c: o_data_a = 16'b1110001100001000;
            14'h306d: o_data_a = 16'b0000000000111101;
            14'h306e: o_data_a = 16'b1110110000010000;
            14'h306f: o_data_a = 16'b0000000000000000;
            14'h3070: o_data_a = 16'b1111110111101000;
            14'h3071: o_data_a = 16'b1110110010100000;
            14'h3072: o_data_a = 16'b1110001100001000;
            14'h3073: o_data_a = 16'b0000000000000000;
            14'h3074: o_data_a = 16'b1111110111001000;
            14'h3075: o_data_a = 16'b1111110010100000;
            14'h3076: o_data_a = 16'b1110101010001000;
            14'h3077: o_data_a = 16'b0000000000000000;
            14'h3078: o_data_a = 16'b1111110111001000;
            14'h3079: o_data_a = 16'b1111110010100000;
            14'h307a: o_data_a = 16'b1110101010001000;
            14'h307b: o_data_a = 16'b0000000000000000;
            14'h307c: o_data_a = 16'b1111110111001000;
            14'h307d: o_data_a = 16'b1111110010100000;
            14'h307e: o_data_a = 16'b1110101010001000;
            14'h307f: o_data_a = 16'b0000000000111111;
            14'h3080: o_data_a = 16'b1110110000010000;
            14'h3081: o_data_a = 16'b0000000000000000;
            14'h3082: o_data_a = 16'b1111110111101000;
            14'h3083: o_data_a = 16'b1110110010100000;
            14'h3084: o_data_a = 16'b1110001100001000;
            14'h3085: o_data_a = 16'b0000000000000000;
            14'h3086: o_data_a = 16'b1111110111001000;
            14'h3087: o_data_a = 16'b1111110010100000;
            14'h3088: o_data_a = 16'b1110101010001000;
            14'h3089: o_data_a = 16'b0000000000000000;
            14'h308a: o_data_a = 16'b1111110111001000;
            14'h308b: o_data_a = 16'b1111110010100000;
            14'h308c: o_data_a = 16'b1110101010001000;
            14'h308d: o_data_a = 16'b0000000000111111;
            14'h308e: o_data_a = 16'b1110110000010000;
            14'h308f: o_data_a = 16'b0000000000000000;
            14'h3090: o_data_a = 16'b1111110111101000;
            14'h3091: o_data_a = 16'b1110110010100000;
            14'h3092: o_data_a = 16'b1110001100001000;
            14'h3093: o_data_a = 16'b0000000000000000;
            14'h3094: o_data_a = 16'b1111110111001000;
            14'h3095: o_data_a = 16'b1111110010100000;
            14'h3096: o_data_a = 16'b1110101010001000;
            14'h3097: o_data_a = 16'b0000000000000000;
            14'h3098: o_data_a = 16'b1111110111001000;
            14'h3099: o_data_a = 16'b1111110010100000;
            14'h309a: o_data_a = 16'b1110101010001000;
            14'h309b: o_data_a = 16'b0000000000000000;
            14'h309c: o_data_a = 16'b1111110111001000;
            14'h309d: o_data_a = 16'b1111110010100000;
            14'h309e: o_data_a = 16'b1110101010001000;
            14'h309f: o_data_a = 16'b0000000000000000;
            14'h30a0: o_data_a = 16'b1111110111001000;
            14'h30a1: o_data_a = 16'b1111110010100000;
            14'h30a2: o_data_a = 16'b1110101010001000;
            14'h30a3: o_data_a = 16'b0000000000001100;
            14'h30a4: o_data_a = 16'b1110110000010000;
            14'h30a5: o_data_a = 16'b0000000000001101;
            14'h30a6: o_data_a = 16'b1110001100001000;
            14'h30a7: o_data_a = 16'b0100010110110011;
            14'h30a8: o_data_a = 16'b1110110000010000;
            14'h30a9: o_data_a = 16'b0000000000001110;
            14'h30aa: o_data_a = 16'b1110001100001000;
            14'h30ab: o_data_a = 16'b0011000010101111;
            14'h30ac: o_data_a = 16'b1110110000010000;
            14'h30ad: o_data_a = 16'b0000000001011111;
            14'h30ae: o_data_a = 16'b1110101010000111;
            14'h30af: o_data_a = 16'b0000000000000000;
            14'h30b0: o_data_a = 16'b1111110010101000;
            14'h30b1: o_data_a = 16'b1111110000010000;
            14'h30b2: o_data_a = 16'b0000000000000101;
            14'h30b3: o_data_a = 16'b1110001100001000;
            14'h30b4: o_data_a = 16'b0000000000111110;
            14'h30b5: o_data_a = 16'b1110110000010000;
            14'h30b6: o_data_a = 16'b0000000000000000;
            14'h30b7: o_data_a = 16'b1111110111101000;
            14'h30b8: o_data_a = 16'b1110110010100000;
            14'h30b9: o_data_a = 16'b1110001100001000;
            14'h30ba: o_data_a = 16'b0000000000000000;
            14'h30bb: o_data_a = 16'b1111110111001000;
            14'h30bc: o_data_a = 16'b1111110010100000;
            14'h30bd: o_data_a = 16'b1110101010001000;
            14'h30be: o_data_a = 16'b0000000000000000;
            14'h30bf: o_data_a = 16'b1111110111001000;
            14'h30c0: o_data_a = 16'b1111110010100000;
            14'h30c1: o_data_a = 16'b1110101010001000;
            14'h30c2: o_data_a = 16'b0000000000000011;
            14'h30c3: o_data_a = 16'b1110110000010000;
            14'h30c4: o_data_a = 16'b0000000000000000;
            14'h30c5: o_data_a = 16'b1111110111101000;
            14'h30c6: o_data_a = 16'b1110110010100000;
            14'h30c7: o_data_a = 16'b1110001100001000;
            14'h30c8: o_data_a = 16'b0000000000000110;
            14'h30c9: o_data_a = 16'b1110110000010000;
            14'h30ca: o_data_a = 16'b0000000000000000;
            14'h30cb: o_data_a = 16'b1111110111101000;
            14'h30cc: o_data_a = 16'b1110110010100000;
            14'h30cd: o_data_a = 16'b1110001100001000;
            14'h30ce: o_data_a = 16'b0000000000001100;
            14'h30cf: o_data_a = 16'b1110110000010000;
            14'h30d0: o_data_a = 16'b0000000000000000;
            14'h30d1: o_data_a = 16'b1111110111101000;
            14'h30d2: o_data_a = 16'b1110110010100000;
            14'h30d3: o_data_a = 16'b1110001100001000;
            14'h30d4: o_data_a = 16'b0000000000011000;
            14'h30d5: o_data_a = 16'b1110110000010000;
            14'h30d6: o_data_a = 16'b0000000000000000;
            14'h30d7: o_data_a = 16'b1111110111101000;
            14'h30d8: o_data_a = 16'b1110110010100000;
            14'h30d9: o_data_a = 16'b1110001100001000;
            14'h30da: o_data_a = 16'b0000000000001100;
            14'h30db: o_data_a = 16'b1110110000010000;
            14'h30dc: o_data_a = 16'b0000000000000000;
            14'h30dd: o_data_a = 16'b1111110111101000;
            14'h30de: o_data_a = 16'b1110110010100000;
            14'h30df: o_data_a = 16'b1110001100001000;
            14'h30e0: o_data_a = 16'b0000000000000110;
            14'h30e1: o_data_a = 16'b1110110000010000;
            14'h30e2: o_data_a = 16'b0000000000000000;
            14'h30e3: o_data_a = 16'b1111110111101000;
            14'h30e4: o_data_a = 16'b1110110010100000;
            14'h30e5: o_data_a = 16'b1110001100001000;
            14'h30e6: o_data_a = 16'b0000000000000011;
            14'h30e7: o_data_a = 16'b1110110000010000;
            14'h30e8: o_data_a = 16'b0000000000000000;
            14'h30e9: o_data_a = 16'b1111110111101000;
            14'h30ea: o_data_a = 16'b1110110010100000;
            14'h30eb: o_data_a = 16'b1110001100001000;
            14'h30ec: o_data_a = 16'b0000000000000000;
            14'h30ed: o_data_a = 16'b1111110111001000;
            14'h30ee: o_data_a = 16'b1111110010100000;
            14'h30ef: o_data_a = 16'b1110101010001000;
            14'h30f0: o_data_a = 16'b0000000000000000;
            14'h30f1: o_data_a = 16'b1111110111001000;
            14'h30f2: o_data_a = 16'b1111110010100000;
            14'h30f3: o_data_a = 16'b1110101010001000;
            14'h30f4: o_data_a = 16'b0000000000001100;
            14'h30f5: o_data_a = 16'b1110110000010000;
            14'h30f6: o_data_a = 16'b0000000000001101;
            14'h30f7: o_data_a = 16'b1110001100001000;
            14'h30f8: o_data_a = 16'b0100010110110011;
            14'h30f9: o_data_a = 16'b1110110000010000;
            14'h30fa: o_data_a = 16'b0000000000001110;
            14'h30fb: o_data_a = 16'b1110001100001000;
            14'h30fc: o_data_a = 16'b0011000100000000;
            14'h30fd: o_data_a = 16'b1110110000010000;
            14'h30fe: o_data_a = 16'b0000000001011111;
            14'h30ff: o_data_a = 16'b1110101010000111;
            14'h3100: o_data_a = 16'b0000000000000000;
            14'h3101: o_data_a = 16'b1111110010101000;
            14'h3102: o_data_a = 16'b1111110000010000;
            14'h3103: o_data_a = 16'b0000000000000101;
            14'h3104: o_data_a = 16'b1110001100001000;
            14'h3105: o_data_a = 16'b0000000001000000;
            14'h3106: o_data_a = 16'b1110110000010000;
            14'h3107: o_data_a = 16'b0000000000000000;
            14'h3108: o_data_a = 16'b1111110111101000;
            14'h3109: o_data_a = 16'b1110110010100000;
            14'h310a: o_data_a = 16'b1110001100001000;
            14'h310b: o_data_a = 16'b0000000000011110;
            14'h310c: o_data_a = 16'b1110110000010000;
            14'h310d: o_data_a = 16'b0000000000000000;
            14'h310e: o_data_a = 16'b1111110111101000;
            14'h310f: o_data_a = 16'b1110110010100000;
            14'h3110: o_data_a = 16'b1110001100001000;
            14'h3111: o_data_a = 16'b0000000000110011;
            14'h3112: o_data_a = 16'b1110110000010000;
            14'h3113: o_data_a = 16'b0000000000000000;
            14'h3114: o_data_a = 16'b1111110111101000;
            14'h3115: o_data_a = 16'b1110110010100000;
            14'h3116: o_data_a = 16'b1110001100001000;
            14'h3117: o_data_a = 16'b0000000000110011;
            14'h3118: o_data_a = 16'b1110110000010000;
            14'h3119: o_data_a = 16'b0000000000000000;
            14'h311a: o_data_a = 16'b1111110111101000;
            14'h311b: o_data_a = 16'b1110110010100000;
            14'h311c: o_data_a = 16'b1110001100001000;
            14'h311d: o_data_a = 16'b0000000000111011;
            14'h311e: o_data_a = 16'b1110110000010000;
            14'h311f: o_data_a = 16'b0000000000000000;
            14'h3120: o_data_a = 16'b1111110111101000;
            14'h3121: o_data_a = 16'b1110110010100000;
            14'h3122: o_data_a = 16'b1110001100001000;
            14'h3123: o_data_a = 16'b0000000000111011;
            14'h3124: o_data_a = 16'b1110110000010000;
            14'h3125: o_data_a = 16'b0000000000000000;
            14'h3126: o_data_a = 16'b1111110111101000;
            14'h3127: o_data_a = 16'b1110110010100000;
            14'h3128: o_data_a = 16'b1110001100001000;
            14'h3129: o_data_a = 16'b0000000000111011;
            14'h312a: o_data_a = 16'b1110110000010000;
            14'h312b: o_data_a = 16'b0000000000000000;
            14'h312c: o_data_a = 16'b1111110111101000;
            14'h312d: o_data_a = 16'b1110110010100000;
            14'h312e: o_data_a = 16'b1110001100001000;
            14'h312f: o_data_a = 16'b0000000000011011;
            14'h3130: o_data_a = 16'b1110110000010000;
            14'h3131: o_data_a = 16'b0000000000000000;
            14'h3132: o_data_a = 16'b1111110111101000;
            14'h3133: o_data_a = 16'b1110110010100000;
            14'h3134: o_data_a = 16'b1110001100001000;
            14'h3135: o_data_a = 16'b0000000000000011;
            14'h3136: o_data_a = 16'b1110110000010000;
            14'h3137: o_data_a = 16'b0000000000000000;
            14'h3138: o_data_a = 16'b1111110111101000;
            14'h3139: o_data_a = 16'b1110110010100000;
            14'h313a: o_data_a = 16'b1110001100001000;
            14'h313b: o_data_a = 16'b0000000000011110;
            14'h313c: o_data_a = 16'b1110110000010000;
            14'h313d: o_data_a = 16'b0000000000000000;
            14'h313e: o_data_a = 16'b1111110111101000;
            14'h313f: o_data_a = 16'b1110110010100000;
            14'h3140: o_data_a = 16'b1110001100001000;
            14'h3141: o_data_a = 16'b0000000000000000;
            14'h3142: o_data_a = 16'b1111110111001000;
            14'h3143: o_data_a = 16'b1111110010100000;
            14'h3144: o_data_a = 16'b1110101010001000;
            14'h3145: o_data_a = 16'b0000000000000000;
            14'h3146: o_data_a = 16'b1111110111001000;
            14'h3147: o_data_a = 16'b1111110010100000;
            14'h3148: o_data_a = 16'b1110101010001000;
            14'h3149: o_data_a = 16'b0000000000001100;
            14'h314a: o_data_a = 16'b1110110000010000;
            14'h314b: o_data_a = 16'b0000000000001101;
            14'h314c: o_data_a = 16'b1110001100001000;
            14'h314d: o_data_a = 16'b0100010110110011;
            14'h314e: o_data_a = 16'b1110110000010000;
            14'h314f: o_data_a = 16'b0000000000001110;
            14'h3150: o_data_a = 16'b1110001100001000;
            14'h3151: o_data_a = 16'b0011000101010101;
            14'h3152: o_data_a = 16'b1110110000010000;
            14'h3153: o_data_a = 16'b0000000001011111;
            14'h3154: o_data_a = 16'b1110101010000111;
            14'h3155: o_data_a = 16'b0000000000000000;
            14'h3156: o_data_a = 16'b1111110010101000;
            14'h3157: o_data_a = 16'b1111110000010000;
            14'h3158: o_data_a = 16'b0000000000000101;
            14'h3159: o_data_a = 16'b1110001100001000;
            14'h315a: o_data_a = 16'b0000000000111111;
            14'h315b: o_data_a = 16'b1110110000010000;
            14'h315c: o_data_a = 16'b0000000000000000;
            14'h315d: o_data_a = 16'b1111110111101000;
            14'h315e: o_data_a = 16'b1110110010100000;
            14'h315f: o_data_a = 16'b1110001100001000;
            14'h3160: o_data_a = 16'b0000000000011110;
            14'h3161: o_data_a = 16'b1110110000010000;
            14'h3162: o_data_a = 16'b0000000000000000;
            14'h3163: o_data_a = 16'b1111110111101000;
            14'h3164: o_data_a = 16'b1110110010100000;
            14'h3165: o_data_a = 16'b1110001100001000;
            14'h3166: o_data_a = 16'b0000000000110011;
            14'h3167: o_data_a = 16'b1110110000010000;
            14'h3168: o_data_a = 16'b0000000000000000;
            14'h3169: o_data_a = 16'b1111110111101000;
            14'h316a: o_data_a = 16'b1110110010100000;
            14'h316b: o_data_a = 16'b1110001100001000;
            14'h316c: o_data_a = 16'b0000000000110011;
            14'h316d: o_data_a = 16'b1110110000010000;
            14'h316e: o_data_a = 16'b0000000000000000;
            14'h316f: o_data_a = 16'b1111110111101000;
            14'h3170: o_data_a = 16'b1110110010100000;
            14'h3171: o_data_a = 16'b1110001100001000;
            14'h3172: o_data_a = 16'b0000000000011000;
            14'h3173: o_data_a = 16'b1110110000010000;
            14'h3174: o_data_a = 16'b0000000000000000;
            14'h3175: o_data_a = 16'b1111110111101000;
            14'h3176: o_data_a = 16'b1110110010100000;
            14'h3177: o_data_a = 16'b1110001100001000;
            14'h3178: o_data_a = 16'b0000000000001100;
            14'h3179: o_data_a = 16'b1110110000010000;
            14'h317a: o_data_a = 16'b0000000000000000;
            14'h317b: o_data_a = 16'b1111110111101000;
            14'h317c: o_data_a = 16'b1110110010100000;
            14'h317d: o_data_a = 16'b1110001100001000;
            14'h317e: o_data_a = 16'b0000000000001100;
            14'h317f: o_data_a = 16'b1110110000010000;
            14'h3180: o_data_a = 16'b0000000000000000;
            14'h3181: o_data_a = 16'b1111110111101000;
            14'h3182: o_data_a = 16'b1110110010100000;
            14'h3183: o_data_a = 16'b1110001100001000;
            14'h3184: o_data_a = 16'b0000000000000000;
            14'h3185: o_data_a = 16'b1111110111001000;
            14'h3186: o_data_a = 16'b1111110010100000;
            14'h3187: o_data_a = 16'b1110101010001000;
            14'h3188: o_data_a = 16'b0000000000001100;
            14'h3189: o_data_a = 16'b1110110000010000;
            14'h318a: o_data_a = 16'b0000000000000000;
            14'h318b: o_data_a = 16'b1111110111101000;
            14'h318c: o_data_a = 16'b1110110010100000;
            14'h318d: o_data_a = 16'b1110001100001000;
            14'h318e: o_data_a = 16'b0000000000001100;
            14'h318f: o_data_a = 16'b1110110000010000;
            14'h3190: o_data_a = 16'b0000000000000000;
            14'h3191: o_data_a = 16'b1111110111101000;
            14'h3192: o_data_a = 16'b1110110010100000;
            14'h3193: o_data_a = 16'b1110001100001000;
            14'h3194: o_data_a = 16'b0000000000000000;
            14'h3195: o_data_a = 16'b1111110111001000;
            14'h3196: o_data_a = 16'b1111110010100000;
            14'h3197: o_data_a = 16'b1110101010001000;
            14'h3198: o_data_a = 16'b0000000000000000;
            14'h3199: o_data_a = 16'b1111110111001000;
            14'h319a: o_data_a = 16'b1111110010100000;
            14'h319b: o_data_a = 16'b1110101010001000;
            14'h319c: o_data_a = 16'b0000000000001100;
            14'h319d: o_data_a = 16'b1110110000010000;
            14'h319e: o_data_a = 16'b0000000000001101;
            14'h319f: o_data_a = 16'b1110001100001000;
            14'h31a0: o_data_a = 16'b0100010110110011;
            14'h31a1: o_data_a = 16'b1110110000010000;
            14'h31a2: o_data_a = 16'b0000000000001110;
            14'h31a3: o_data_a = 16'b1110001100001000;
            14'h31a4: o_data_a = 16'b0011000110101000;
            14'h31a5: o_data_a = 16'b1110110000010000;
            14'h31a6: o_data_a = 16'b0000000001011111;
            14'h31a7: o_data_a = 16'b1110101010000111;
            14'h31a8: o_data_a = 16'b0000000000000000;
            14'h31a9: o_data_a = 16'b1111110010101000;
            14'h31aa: o_data_a = 16'b1111110000010000;
            14'h31ab: o_data_a = 16'b0000000000000101;
            14'h31ac: o_data_a = 16'b1110001100001000;
            14'h31ad: o_data_a = 16'b0000000001000001;
            14'h31ae: o_data_a = 16'b1110110000010000;
            14'h31af: o_data_a = 16'b0000000000000000;
            14'h31b0: o_data_a = 16'b1111110111101000;
            14'h31b1: o_data_a = 16'b1110110010100000;
            14'h31b2: o_data_a = 16'b1110001100001000;
            14'h31b3: o_data_a = 16'b0000000000001100;
            14'h31b4: o_data_a = 16'b1110110000010000;
            14'h31b5: o_data_a = 16'b0000000000000000;
            14'h31b6: o_data_a = 16'b1111110111101000;
            14'h31b7: o_data_a = 16'b1110110010100000;
            14'h31b8: o_data_a = 16'b1110001100001000;
            14'h31b9: o_data_a = 16'b0000000000011110;
            14'h31ba: o_data_a = 16'b1110110000010000;
            14'h31bb: o_data_a = 16'b0000000000000000;
            14'h31bc: o_data_a = 16'b1111110111101000;
            14'h31bd: o_data_a = 16'b1110110010100000;
            14'h31be: o_data_a = 16'b1110001100001000;
            14'h31bf: o_data_a = 16'b0000000000110011;
            14'h31c0: o_data_a = 16'b1110110000010000;
            14'h31c1: o_data_a = 16'b0000000000000000;
            14'h31c2: o_data_a = 16'b1111110111101000;
            14'h31c3: o_data_a = 16'b1110110010100000;
            14'h31c4: o_data_a = 16'b1110001100001000;
            14'h31c5: o_data_a = 16'b0000000000110011;
            14'h31c6: o_data_a = 16'b1110110000010000;
            14'h31c7: o_data_a = 16'b0000000000000000;
            14'h31c8: o_data_a = 16'b1111110111101000;
            14'h31c9: o_data_a = 16'b1110110010100000;
            14'h31ca: o_data_a = 16'b1110001100001000;
            14'h31cb: o_data_a = 16'b0000000000111111;
            14'h31cc: o_data_a = 16'b1110110000010000;
            14'h31cd: o_data_a = 16'b0000000000000000;
            14'h31ce: o_data_a = 16'b1111110111101000;
            14'h31cf: o_data_a = 16'b1110110010100000;
            14'h31d0: o_data_a = 16'b1110001100001000;
            14'h31d1: o_data_a = 16'b0000000000110011;
            14'h31d2: o_data_a = 16'b1110110000010000;
            14'h31d3: o_data_a = 16'b0000000000000000;
            14'h31d4: o_data_a = 16'b1111110111101000;
            14'h31d5: o_data_a = 16'b1110110010100000;
            14'h31d6: o_data_a = 16'b1110001100001000;
            14'h31d7: o_data_a = 16'b0000000000110011;
            14'h31d8: o_data_a = 16'b1110110000010000;
            14'h31d9: o_data_a = 16'b0000000000000000;
            14'h31da: o_data_a = 16'b1111110111101000;
            14'h31db: o_data_a = 16'b1110110010100000;
            14'h31dc: o_data_a = 16'b1110001100001000;
            14'h31dd: o_data_a = 16'b0000000000110011;
            14'h31de: o_data_a = 16'b1110110000010000;
            14'h31df: o_data_a = 16'b0000000000000000;
            14'h31e0: o_data_a = 16'b1111110111101000;
            14'h31e1: o_data_a = 16'b1110110010100000;
            14'h31e2: o_data_a = 16'b1110001100001000;
            14'h31e3: o_data_a = 16'b0000000000110011;
            14'h31e4: o_data_a = 16'b1110110000010000;
            14'h31e5: o_data_a = 16'b0000000000000000;
            14'h31e6: o_data_a = 16'b1111110111101000;
            14'h31e7: o_data_a = 16'b1110110010100000;
            14'h31e8: o_data_a = 16'b1110001100001000;
            14'h31e9: o_data_a = 16'b0000000000000000;
            14'h31ea: o_data_a = 16'b1111110111001000;
            14'h31eb: o_data_a = 16'b1111110010100000;
            14'h31ec: o_data_a = 16'b1110101010001000;
            14'h31ed: o_data_a = 16'b0000000000000000;
            14'h31ee: o_data_a = 16'b1111110111001000;
            14'h31ef: o_data_a = 16'b1111110010100000;
            14'h31f0: o_data_a = 16'b1110101010001000;
            14'h31f1: o_data_a = 16'b0000000000001100;
            14'h31f2: o_data_a = 16'b1110110000010000;
            14'h31f3: o_data_a = 16'b0000000000001101;
            14'h31f4: o_data_a = 16'b1110001100001000;
            14'h31f5: o_data_a = 16'b0100010110110011;
            14'h31f6: o_data_a = 16'b1110110000010000;
            14'h31f7: o_data_a = 16'b0000000000001110;
            14'h31f8: o_data_a = 16'b1110001100001000;
            14'h31f9: o_data_a = 16'b0011000111111101;
            14'h31fa: o_data_a = 16'b1110110000010000;
            14'h31fb: o_data_a = 16'b0000000001011111;
            14'h31fc: o_data_a = 16'b1110101010000111;
            14'h31fd: o_data_a = 16'b0000000000000000;
            14'h31fe: o_data_a = 16'b1111110010101000;
            14'h31ff: o_data_a = 16'b1111110000010000;
            14'h3200: o_data_a = 16'b0000000000000101;
            14'h3201: o_data_a = 16'b1110001100001000;
            14'h3202: o_data_a = 16'b0000000001000010;
            14'h3203: o_data_a = 16'b1110110000010000;
            14'h3204: o_data_a = 16'b0000000000000000;
            14'h3205: o_data_a = 16'b1111110111101000;
            14'h3206: o_data_a = 16'b1110110010100000;
            14'h3207: o_data_a = 16'b1110001100001000;
            14'h3208: o_data_a = 16'b0000000000011111;
            14'h3209: o_data_a = 16'b1110110000010000;
            14'h320a: o_data_a = 16'b0000000000000000;
            14'h320b: o_data_a = 16'b1111110111101000;
            14'h320c: o_data_a = 16'b1110110010100000;
            14'h320d: o_data_a = 16'b1110001100001000;
            14'h320e: o_data_a = 16'b0000000000110011;
            14'h320f: o_data_a = 16'b1110110000010000;
            14'h3210: o_data_a = 16'b0000000000000000;
            14'h3211: o_data_a = 16'b1111110111101000;
            14'h3212: o_data_a = 16'b1110110010100000;
            14'h3213: o_data_a = 16'b1110001100001000;
            14'h3214: o_data_a = 16'b0000000000110011;
            14'h3215: o_data_a = 16'b1110110000010000;
            14'h3216: o_data_a = 16'b0000000000000000;
            14'h3217: o_data_a = 16'b1111110111101000;
            14'h3218: o_data_a = 16'b1110110010100000;
            14'h3219: o_data_a = 16'b1110001100001000;
            14'h321a: o_data_a = 16'b0000000000110011;
            14'h321b: o_data_a = 16'b1110110000010000;
            14'h321c: o_data_a = 16'b0000000000000000;
            14'h321d: o_data_a = 16'b1111110111101000;
            14'h321e: o_data_a = 16'b1110110010100000;
            14'h321f: o_data_a = 16'b1110001100001000;
            14'h3220: o_data_a = 16'b0000000000011111;
            14'h3221: o_data_a = 16'b1110110000010000;
            14'h3222: o_data_a = 16'b0000000000000000;
            14'h3223: o_data_a = 16'b1111110111101000;
            14'h3224: o_data_a = 16'b1110110010100000;
            14'h3225: o_data_a = 16'b1110001100001000;
            14'h3226: o_data_a = 16'b0000000000110011;
            14'h3227: o_data_a = 16'b1110110000010000;
            14'h3228: o_data_a = 16'b0000000000000000;
            14'h3229: o_data_a = 16'b1111110111101000;
            14'h322a: o_data_a = 16'b1110110010100000;
            14'h322b: o_data_a = 16'b1110001100001000;
            14'h322c: o_data_a = 16'b0000000000110011;
            14'h322d: o_data_a = 16'b1110110000010000;
            14'h322e: o_data_a = 16'b0000000000000000;
            14'h322f: o_data_a = 16'b1111110111101000;
            14'h3230: o_data_a = 16'b1110110010100000;
            14'h3231: o_data_a = 16'b1110001100001000;
            14'h3232: o_data_a = 16'b0000000000110011;
            14'h3233: o_data_a = 16'b1110110000010000;
            14'h3234: o_data_a = 16'b0000000000000000;
            14'h3235: o_data_a = 16'b1111110111101000;
            14'h3236: o_data_a = 16'b1110110010100000;
            14'h3237: o_data_a = 16'b1110001100001000;
            14'h3238: o_data_a = 16'b0000000000011111;
            14'h3239: o_data_a = 16'b1110110000010000;
            14'h323a: o_data_a = 16'b0000000000000000;
            14'h323b: o_data_a = 16'b1111110111101000;
            14'h323c: o_data_a = 16'b1110110010100000;
            14'h323d: o_data_a = 16'b1110001100001000;
            14'h323e: o_data_a = 16'b0000000000000000;
            14'h323f: o_data_a = 16'b1111110111001000;
            14'h3240: o_data_a = 16'b1111110010100000;
            14'h3241: o_data_a = 16'b1110101010001000;
            14'h3242: o_data_a = 16'b0000000000000000;
            14'h3243: o_data_a = 16'b1111110111001000;
            14'h3244: o_data_a = 16'b1111110010100000;
            14'h3245: o_data_a = 16'b1110101010001000;
            14'h3246: o_data_a = 16'b0000000000001100;
            14'h3247: o_data_a = 16'b1110110000010000;
            14'h3248: o_data_a = 16'b0000000000001101;
            14'h3249: o_data_a = 16'b1110001100001000;
            14'h324a: o_data_a = 16'b0100010110110011;
            14'h324b: o_data_a = 16'b1110110000010000;
            14'h324c: o_data_a = 16'b0000000000001110;
            14'h324d: o_data_a = 16'b1110001100001000;
            14'h324e: o_data_a = 16'b0011001001010010;
            14'h324f: o_data_a = 16'b1110110000010000;
            14'h3250: o_data_a = 16'b0000000001011111;
            14'h3251: o_data_a = 16'b1110101010000111;
            14'h3252: o_data_a = 16'b0000000000000000;
            14'h3253: o_data_a = 16'b1111110010101000;
            14'h3254: o_data_a = 16'b1111110000010000;
            14'h3255: o_data_a = 16'b0000000000000101;
            14'h3256: o_data_a = 16'b1110001100001000;
            14'h3257: o_data_a = 16'b0000000001000011;
            14'h3258: o_data_a = 16'b1110110000010000;
            14'h3259: o_data_a = 16'b0000000000000000;
            14'h325a: o_data_a = 16'b1111110111101000;
            14'h325b: o_data_a = 16'b1110110010100000;
            14'h325c: o_data_a = 16'b1110001100001000;
            14'h325d: o_data_a = 16'b0000000000011100;
            14'h325e: o_data_a = 16'b1110110000010000;
            14'h325f: o_data_a = 16'b0000000000000000;
            14'h3260: o_data_a = 16'b1111110111101000;
            14'h3261: o_data_a = 16'b1110110010100000;
            14'h3262: o_data_a = 16'b1110001100001000;
            14'h3263: o_data_a = 16'b0000000000110110;
            14'h3264: o_data_a = 16'b1110110000010000;
            14'h3265: o_data_a = 16'b0000000000000000;
            14'h3266: o_data_a = 16'b1111110111101000;
            14'h3267: o_data_a = 16'b1110110010100000;
            14'h3268: o_data_a = 16'b1110001100001000;
            14'h3269: o_data_a = 16'b0000000000100011;
            14'h326a: o_data_a = 16'b1110110000010000;
            14'h326b: o_data_a = 16'b0000000000000000;
            14'h326c: o_data_a = 16'b1111110111101000;
            14'h326d: o_data_a = 16'b1110110010100000;
            14'h326e: o_data_a = 16'b1110001100001000;
            14'h326f: o_data_a = 16'b0000000000000011;
            14'h3270: o_data_a = 16'b1110110000010000;
            14'h3271: o_data_a = 16'b0000000000000000;
            14'h3272: o_data_a = 16'b1111110111101000;
            14'h3273: o_data_a = 16'b1110110010100000;
            14'h3274: o_data_a = 16'b1110001100001000;
            14'h3275: o_data_a = 16'b0000000000000011;
            14'h3276: o_data_a = 16'b1110110000010000;
            14'h3277: o_data_a = 16'b0000000000000000;
            14'h3278: o_data_a = 16'b1111110111101000;
            14'h3279: o_data_a = 16'b1110110010100000;
            14'h327a: o_data_a = 16'b1110001100001000;
            14'h327b: o_data_a = 16'b0000000000000011;
            14'h327c: o_data_a = 16'b1110110000010000;
            14'h327d: o_data_a = 16'b0000000000000000;
            14'h327e: o_data_a = 16'b1111110111101000;
            14'h327f: o_data_a = 16'b1110110010100000;
            14'h3280: o_data_a = 16'b1110001100001000;
            14'h3281: o_data_a = 16'b0000000000100011;
            14'h3282: o_data_a = 16'b1110110000010000;
            14'h3283: o_data_a = 16'b0000000000000000;
            14'h3284: o_data_a = 16'b1111110111101000;
            14'h3285: o_data_a = 16'b1110110010100000;
            14'h3286: o_data_a = 16'b1110001100001000;
            14'h3287: o_data_a = 16'b0000000000110110;
            14'h3288: o_data_a = 16'b1110110000010000;
            14'h3289: o_data_a = 16'b0000000000000000;
            14'h328a: o_data_a = 16'b1111110111101000;
            14'h328b: o_data_a = 16'b1110110010100000;
            14'h328c: o_data_a = 16'b1110001100001000;
            14'h328d: o_data_a = 16'b0000000000011100;
            14'h328e: o_data_a = 16'b1110110000010000;
            14'h328f: o_data_a = 16'b0000000000000000;
            14'h3290: o_data_a = 16'b1111110111101000;
            14'h3291: o_data_a = 16'b1110110010100000;
            14'h3292: o_data_a = 16'b1110001100001000;
            14'h3293: o_data_a = 16'b0000000000000000;
            14'h3294: o_data_a = 16'b1111110111001000;
            14'h3295: o_data_a = 16'b1111110010100000;
            14'h3296: o_data_a = 16'b1110101010001000;
            14'h3297: o_data_a = 16'b0000000000000000;
            14'h3298: o_data_a = 16'b1111110111001000;
            14'h3299: o_data_a = 16'b1111110010100000;
            14'h329a: o_data_a = 16'b1110101010001000;
            14'h329b: o_data_a = 16'b0000000000001100;
            14'h329c: o_data_a = 16'b1110110000010000;
            14'h329d: o_data_a = 16'b0000000000001101;
            14'h329e: o_data_a = 16'b1110001100001000;
            14'h329f: o_data_a = 16'b0100010110110011;
            14'h32a0: o_data_a = 16'b1110110000010000;
            14'h32a1: o_data_a = 16'b0000000000001110;
            14'h32a2: o_data_a = 16'b1110001100001000;
            14'h32a3: o_data_a = 16'b0011001010100111;
            14'h32a4: o_data_a = 16'b1110110000010000;
            14'h32a5: o_data_a = 16'b0000000001011111;
            14'h32a6: o_data_a = 16'b1110101010000111;
            14'h32a7: o_data_a = 16'b0000000000000000;
            14'h32a8: o_data_a = 16'b1111110010101000;
            14'h32a9: o_data_a = 16'b1111110000010000;
            14'h32aa: o_data_a = 16'b0000000000000101;
            14'h32ab: o_data_a = 16'b1110001100001000;
            14'h32ac: o_data_a = 16'b0000000001000100;
            14'h32ad: o_data_a = 16'b1110110000010000;
            14'h32ae: o_data_a = 16'b0000000000000000;
            14'h32af: o_data_a = 16'b1111110111101000;
            14'h32b0: o_data_a = 16'b1110110010100000;
            14'h32b1: o_data_a = 16'b1110001100001000;
            14'h32b2: o_data_a = 16'b0000000000001111;
            14'h32b3: o_data_a = 16'b1110110000010000;
            14'h32b4: o_data_a = 16'b0000000000000000;
            14'h32b5: o_data_a = 16'b1111110111101000;
            14'h32b6: o_data_a = 16'b1110110010100000;
            14'h32b7: o_data_a = 16'b1110001100001000;
            14'h32b8: o_data_a = 16'b0000000000011011;
            14'h32b9: o_data_a = 16'b1110110000010000;
            14'h32ba: o_data_a = 16'b0000000000000000;
            14'h32bb: o_data_a = 16'b1111110111101000;
            14'h32bc: o_data_a = 16'b1110110010100000;
            14'h32bd: o_data_a = 16'b1110001100001000;
            14'h32be: o_data_a = 16'b0000000000110011;
            14'h32bf: o_data_a = 16'b1110110000010000;
            14'h32c0: o_data_a = 16'b0000000000000000;
            14'h32c1: o_data_a = 16'b1111110111101000;
            14'h32c2: o_data_a = 16'b1110110010100000;
            14'h32c3: o_data_a = 16'b1110001100001000;
            14'h32c4: o_data_a = 16'b0000000000110011;
            14'h32c5: o_data_a = 16'b1110110000010000;
            14'h32c6: o_data_a = 16'b0000000000000000;
            14'h32c7: o_data_a = 16'b1111110111101000;
            14'h32c8: o_data_a = 16'b1110110010100000;
            14'h32c9: o_data_a = 16'b1110001100001000;
            14'h32ca: o_data_a = 16'b0000000000110011;
            14'h32cb: o_data_a = 16'b1110110000010000;
            14'h32cc: o_data_a = 16'b0000000000000000;
            14'h32cd: o_data_a = 16'b1111110111101000;
            14'h32ce: o_data_a = 16'b1110110010100000;
            14'h32cf: o_data_a = 16'b1110001100001000;
            14'h32d0: o_data_a = 16'b0000000000110011;
            14'h32d1: o_data_a = 16'b1110110000010000;
            14'h32d2: o_data_a = 16'b0000000000000000;
            14'h32d3: o_data_a = 16'b1111110111101000;
            14'h32d4: o_data_a = 16'b1110110010100000;
            14'h32d5: o_data_a = 16'b1110001100001000;
            14'h32d6: o_data_a = 16'b0000000000110011;
            14'h32d7: o_data_a = 16'b1110110000010000;
            14'h32d8: o_data_a = 16'b0000000000000000;
            14'h32d9: o_data_a = 16'b1111110111101000;
            14'h32da: o_data_a = 16'b1110110010100000;
            14'h32db: o_data_a = 16'b1110001100001000;
            14'h32dc: o_data_a = 16'b0000000000011011;
            14'h32dd: o_data_a = 16'b1110110000010000;
            14'h32de: o_data_a = 16'b0000000000000000;
            14'h32df: o_data_a = 16'b1111110111101000;
            14'h32e0: o_data_a = 16'b1110110010100000;
            14'h32e1: o_data_a = 16'b1110001100001000;
            14'h32e2: o_data_a = 16'b0000000000001111;
            14'h32e3: o_data_a = 16'b1110110000010000;
            14'h32e4: o_data_a = 16'b0000000000000000;
            14'h32e5: o_data_a = 16'b1111110111101000;
            14'h32e6: o_data_a = 16'b1110110010100000;
            14'h32e7: o_data_a = 16'b1110001100001000;
            14'h32e8: o_data_a = 16'b0000000000000000;
            14'h32e9: o_data_a = 16'b1111110111001000;
            14'h32ea: o_data_a = 16'b1111110010100000;
            14'h32eb: o_data_a = 16'b1110101010001000;
            14'h32ec: o_data_a = 16'b0000000000000000;
            14'h32ed: o_data_a = 16'b1111110111001000;
            14'h32ee: o_data_a = 16'b1111110010100000;
            14'h32ef: o_data_a = 16'b1110101010001000;
            14'h32f0: o_data_a = 16'b0000000000001100;
            14'h32f1: o_data_a = 16'b1110110000010000;
            14'h32f2: o_data_a = 16'b0000000000001101;
            14'h32f3: o_data_a = 16'b1110001100001000;
            14'h32f4: o_data_a = 16'b0100010110110011;
            14'h32f5: o_data_a = 16'b1110110000010000;
            14'h32f6: o_data_a = 16'b0000000000001110;
            14'h32f7: o_data_a = 16'b1110001100001000;
            14'h32f8: o_data_a = 16'b0011001011111100;
            14'h32f9: o_data_a = 16'b1110110000010000;
            14'h32fa: o_data_a = 16'b0000000001011111;
            14'h32fb: o_data_a = 16'b1110101010000111;
            14'h32fc: o_data_a = 16'b0000000000000000;
            14'h32fd: o_data_a = 16'b1111110010101000;
            14'h32fe: o_data_a = 16'b1111110000010000;
            14'h32ff: o_data_a = 16'b0000000000000101;
            14'h3300: o_data_a = 16'b1110001100001000;
            14'h3301: o_data_a = 16'b0000000001000101;
            14'h3302: o_data_a = 16'b1110110000010000;
            14'h3303: o_data_a = 16'b0000000000000000;
            14'h3304: o_data_a = 16'b1111110111101000;
            14'h3305: o_data_a = 16'b1110110010100000;
            14'h3306: o_data_a = 16'b1110001100001000;
            14'h3307: o_data_a = 16'b0000000000111111;
            14'h3308: o_data_a = 16'b1110110000010000;
            14'h3309: o_data_a = 16'b0000000000000000;
            14'h330a: o_data_a = 16'b1111110111101000;
            14'h330b: o_data_a = 16'b1110110010100000;
            14'h330c: o_data_a = 16'b1110001100001000;
            14'h330d: o_data_a = 16'b0000000000110011;
            14'h330e: o_data_a = 16'b1110110000010000;
            14'h330f: o_data_a = 16'b0000000000000000;
            14'h3310: o_data_a = 16'b1111110111101000;
            14'h3311: o_data_a = 16'b1110110010100000;
            14'h3312: o_data_a = 16'b1110001100001000;
            14'h3313: o_data_a = 16'b0000000000100011;
            14'h3314: o_data_a = 16'b1110110000010000;
            14'h3315: o_data_a = 16'b0000000000000000;
            14'h3316: o_data_a = 16'b1111110111101000;
            14'h3317: o_data_a = 16'b1110110010100000;
            14'h3318: o_data_a = 16'b1110001100001000;
            14'h3319: o_data_a = 16'b0000000000001011;
            14'h331a: o_data_a = 16'b1110110000010000;
            14'h331b: o_data_a = 16'b0000000000000000;
            14'h331c: o_data_a = 16'b1111110111101000;
            14'h331d: o_data_a = 16'b1110110010100000;
            14'h331e: o_data_a = 16'b1110001100001000;
            14'h331f: o_data_a = 16'b0000000000001111;
            14'h3320: o_data_a = 16'b1110110000010000;
            14'h3321: o_data_a = 16'b0000000000000000;
            14'h3322: o_data_a = 16'b1111110111101000;
            14'h3323: o_data_a = 16'b1110110010100000;
            14'h3324: o_data_a = 16'b1110001100001000;
            14'h3325: o_data_a = 16'b0000000000001011;
            14'h3326: o_data_a = 16'b1110110000010000;
            14'h3327: o_data_a = 16'b0000000000000000;
            14'h3328: o_data_a = 16'b1111110111101000;
            14'h3329: o_data_a = 16'b1110110010100000;
            14'h332a: o_data_a = 16'b1110001100001000;
            14'h332b: o_data_a = 16'b0000000000100011;
            14'h332c: o_data_a = 16'b1110110000010000;
            14'h332d: o_data_a = 16'b0000000000000000;
            14'h332e: o_data_a = 16'b1111110111101000;
            14'h332f: o_data_a = 16'b1110110010100000;
            14'h3330: o_data_a = 16'b1110001100001000;
            14'h3331: o_data_a = 16'b0000000000110011;
            14'h3332: o_data_a = 16'b1110110000010000;
            14'h3333: o_data_a = 16'b0000000000000000;
            14'h3334: o_data_a = 16'b1111110111101000;
            14'h3335: o_data_a = 16'b1110110010100000;
            14'h3336: o_data_a = 16'b1110001100001000;
            14'h3337: o_data_a = 16'b0000000000111111;
            14'h3338: o_data_a = 16'b1110110000010000;
            14'h3339: o_data_a = 16'b0000000000000000;
            14'h333a: o_data_a = 16'b1111110111101000;
            14'h333b: o_data_a = 16'b1110110010100000;
            14'h333c: o_data_a = 16'b1110001100001000;
            14'h333d: o_data_a = 16'b0000000000000000;
            14'h333e: o_data_a = 16'b1111110111001000;
            14'h333f: o_data_a = 16'b1111110010100000;
            14'h3340: o_data_a = 16'b1110101010001000;
            14'h3341: o_data_a = 16'b0000000000000000;
            14'h3342: o_data_a = 16'b1111110111001000;
            14'h3343: o_data_a = 16'b1111110010100000;
            14'h3344: o_data_a = 16'b1110101010001000;
            14'h3345: o_data_a = 16'b0000000000001100;
            14'h3346: o_data_a = 16'b1110110000010000;
            14'h3347: o_data_a = 16'b0000000000001101;
            14'h3348: o_data_a = 16'b1110001100001000;
            14'h3349: o_data_a = 16'b0100010110110011;
            14'h334a: o_data_a = 16'b1110110000010000;
            14'h334b: o_data_a = 16'b0000000000001110;
            14'h334c: o_data_a = 16'b1110001100001000;
            14'h334d: o_data_a = 16'b0011001101010001;
            14'h334e: o_data_a = 16'b1110110000010000;
            14'h334f: o_data_a = 16'b0000000001011111;
            14'h3350: o_data_a = 16'b1110101010000111;
            14'h3351: o_data_a = 16'b0000000000000000;
            14'h3352: o_data_a = 16'b1111110010101000;
            14'h3353: o_data_a = 16'b1111110000010000;
            14'h3354: o_data_a = 16'b0000000000000101;
            14'h3355: o_data_a = 16'b1110001100001000;
            14'h3356: o_data_a = 16'b0000000001000110;
            14'h3357: o_data_a = 16'b1110110000010000;
            14'h3358: o_data_a = 16'b0000000000000000;
            14'h3359: o_data_a = 16'b1111110111101000;
            14'h335a: o_data_a = 16'b1110110010100000;
            14'h335b: o_data_a = 16'b1110001100001000;
            14'h335c: o_data_a = 16'b0000000000111111;
            14'h335d: o_data_a = 16'b1110110000010000;
            14'h335e: o_data_a = 16'b0000000000000000;
            14'h335f: o_data_a = 16'b1111110111101000;
            14'h3360: o_data_a = 16'b1110110010100000;
            14'h3361: o_data_a = 16'b1110001100001000;
            14'h3362: o_data_a = 16'b0000000000110011;
            14'h3363: o_data_a = 16'b1110110000010000;
            14'h3364: o_data_a = 16'b0000000000000000;
            14'h3365: o_data_a = 16'b1111110111101000;
            14'h3366: o_data_a = 16'b1110110010100000;
            14'h3367: o_data_a = 16'b1110001100001000;
            14'h3368: o_data_a = 16'b0000000000100011;
            14'h3369: o_data_a = 16'b1110110000010000;
            14'h336a: o_data_a = 16'b0000000000000000;
            14'h336b: o_data_a = 16'b1111110111101000;
            14'h336c: o_data_a = 16'b1110110010100000;
            14'h336d: o_data_a = 16'b1110001100001000;
            14'h336e: o_data_a = 16'b0000000000001011;
            14'h336f: o_data_a = 16'b1110110000010000;
            14'h3370: o_data_a = 16'b0000000000000000;
            14'h3371: o_data_a = 16'b1111110111101000;
            14'h3372: o_data_a = 16'b1110110010100000;
            14'h3373: o_data_a = 16'b1110001100001000;
            14'h3374: o_data_a = 16'b0000000000001111;
            14'h3375: o_data_a = 16'b1110110000010000;
            14'h3376: o_data_a = 16'b0000000000000000;
            14'h3377: o_data_a = 16'b1111110111101000;
            14'h3378: o_data_a = 16'b1110110010100000;
            14'h3379: o_data_a = 16'b1110001100001000;
            14'h337a: o_data_a = 16'b0000000000001011;
            14'h337b: o_data_a = 16'b1110110000010000;
            14'h337c: o_data_a = 16'b0000000000000000;
            14'h337d: o_data_a = 16'b1111110111101000;
            14'h337e: o_data_a = 16'b1110110010100000;
            14'h337f: o_data_a = 16'b1110001100001000;
            14'h3380: o_data_a = 16'b0000000000000011;
            14'h3381: o_data_a = 16'b1110110000010000;
            14'h3382: o_data_a = 16'b0000000000000000;
            14'h3383: o_data_a = 16'b1111110111101000;
            14'h3384: o_data_a = 16'b1110110010100000;
            14'h3385: o_data_a = 16'b1110001100001000;
            14'h3386: o_data_a = 16'b0000000000000011;
            14'h3387: o_data_a = 16'b1110110000010000;
            14'h3388: o_data_a = 16'b0000000000000000;
            14'h3389: o_data_a = 16'b1111110111101000;
            14'h338a: o_data_a = 16'b1110110010100000;
            14'h338b: o_data_a = 16'b1110001100001000;
            14'h338c: o_data_a = 16'b0000000000000011;
            14'h338d: o_data_a = 16'b1110110000010000;
            14'h338e: o_data_a = 16'b0000000000000000;
            14'h338f: o_data_a = 16'b1111110111101000;
            14'h3390: o_data_a = 16'b1110110010100000;
            14'h3391: o_data_a = 16'b1110001100001000;
            14'h3392: o_data_a = 16'b0000000000000000;
            14'h3393: o_data_a = 16'b1111110111001000;
            14'h3394: o_data_a = 16'b1111110010100000;
            14'h3395: o_data_a = 16'b1110101010001000;
            14'h3396: o_data_a = 16'b0000000000000000;
            14'h3397: o_data_a = 16'b1111110111001000;
            14'h3398: o_data_a = 16'b1111110010100000;
            14'h3399: o_data_a = 16'b1110101010001000;
            14'h339a: o_data_a = 16'b0000000000001100;
            14'h339b: o_data_a = 16'b1110110000010000;
            14'h339c: o_data_a = 16'b0000000000001101;
            14'h339d: o_data_a = 16'b1110001100001000;
            14'h339e: o_data_a = 16'b0100010110110011;
            14'h339f: o_data_a = 16'b1110110000010000;
            14'h33a0: o_data_a = 16'b0000000000001110;
            14'h33a1: o_data_a = 16'b1110001100001000;
            14'h33a2: o_data_a = 16'b0011001110100110;
            14'h33a3: o_data_a = 16'b1110110000010000;
            14'h33a4: o_data_a = 16'b0000000001011111;
            14'h33a5: o_data_a = 16'b1110101010000111;
            14'h33a6: o_data_a = 16'b0000000000000000;
            14'h33a7: o_data_a = 16'b1111110010101000;
            14'h33a8: o_data_a = 16'b1111110000010000;
            14'h33a9: o_data_a = 16'b0000000000000101;
            14'h33aa: o_data_a = 16'b1110001100001000;
            14'h33ab: o_data_a = 16'b0000000001000111;
            14'h33ac: o_data_a = 16'b1110110000010000;
            14'h33ad: o_data_a = 16'b0000000000000000;
            14'h33ae: o_data_a = 16'b1111110111101000;
            14'h33af: o_data_a = 16'b1110110010100000;
            14'h33b0: o_data_a = 16'b1110001100001000;
            14'h33b1: o_data_a = 16'b0000000000011100;
            14'h33b2: o_data_a = 16'b1110110000010000;
            14'h33b3: o_data_a = 16'b0000000000000000;
            14'h33b4: o_data_a = 16'b1111110111101000;
            14'h33b5: o_data_a = 16'b1110110010100000;
            14'h33b6: o_data_a = 16'b1110001100001000;
            14'h33b7: o_data_a = 16'b0000000000110110;
            14'h33b8: o_data_a = 16'b1110110000010000;
            14'h33b9: o_data_a = 16'b0000000000000000;
            14'h33ba: o_data_a = 16'b1111110111101000;
            14'h33bb: o_data_a = 16'b1110110010100000;
            14'h33bc: o_data_a = 16'b1110001100001000;
            14'h33bd: o_data_a = 16'b0000000000100011;
            14'h33be: o_data_a = 16'b1110110000010000;
            14'h33bf: o_data_a = 16'b0000000000000000;
            14'h33c0: o_data_a = 16'b1111110111101000;
            14'h33c1: o_data_a = 16'b1110110010100000;
            14'h33c2: o_data_a = 16'b1110001100001000;
            14'h33c3: o_data_a = 16'b0000000000000011;
            14'h33c4: o_data_a = 16'b1110110000010000;
            14'h33c5: o_data_a = 16'b0000000000000000;
            14'h33c6: o_data_a = 16'b1111110111101000;
            14'h33c7: o_data_a = 16'b1110110010100000;
            14'h33c8: o_data_a = 16'b1110001100001000;
            14'h33c9: o_data_a = 16'b0000000000111011;
            14'h33ca: o_data_a = 16'b1110110000010000;
            14'h33cb: o_data_a = 16'b0000000000000000;
            14'h33cc: o_data_a = 16'b1111110111101000;
            14'h33cd: o_data_a = 16'b1110110010100000;
            14'h33ce: o_data_a = 16'b1110001100001000;
            14'h33cf: o_data_a = 16'b0000000000110011;
            14'h33d0: o_data_a = 16'b1110110000010000;
            14'h33d1: o_data_a = 16'b0000000000000000;
            14'h33d2: o_data_a = 16'b1111110111101000;
            14'h33d3: o_data_a = 16'b1110110010100000;
            14'h33d4: o_data_a = 16'b1110001100001000;
            14'h33d5: o_data_a = 16'b0000000000110011;
            14'h33d6: o_data_a = 16'b1110110000010000;
            14'h33d7: o_data_a = 16'b0000000000000000;
            14'h33d8: o_data_a = 16'b1111110111101000;
            14'h33d9: o_data_a = 16'b1110110010100000;
            14'h33da: o_data_a = 16'b1110001100001000;
            14'h33db: o_data_a = 16'b0000000000110110;
            14'h33dc: o_data_a = 16'b1110110000010000;
            14'h33dd: o_data_a = 16'b0000000000000000;
            14'h33de: o_data_a = 16'b1111110111101000;
            14'h33df: o_data_a = 16'b1110110010100000;
            14'h33e0: o_data_a = 16'b1110001100001000;
            14'h33e1: o_data_a = 16'b0000000000101100;
            14'h33e2: o_data_a = 16'b1110110000010000;
            14'h33e3: o_data_a = 16'b0000000000000000;
            14'h33e4: o_data_a = 16'b1111110111101000;
            14'h33e5: o_data_a = 16'b1110110010100000;
            14'h33e6: o_data_a = 16'b1110001100001000;
            14'h33e7: o_data_a = 16'b0000000000000000;
            14'h33e8: o_data_a = 16'b1111110111001000;
            14'h33e9: o_data_a = 16'b1111110010100000;
            14'h33ea: o_data_a = 16'b1110101010001000;
            14'h33eb: o_data_a = 16'b0000000000000000;
            14'h33ec: o_data_a = 16'b1111110111001000;
            14'h33ed: o_data_a = 16'b1111110010100000;
            14'h33ee: o_data_a = 16'b1110101010001000;
            14'h33ef: o_data_a = 16'b0000000000001100;
            14'h33f0: o_data_a = 16'b1110110000010000;
            14'h33f1: o_data_a = 16'b0000000000001101;
            14'h33f2: o_data_a = 16'b1110001100001000;
            14'h33f3: o_data_a = 16'b0100010110110011;
            14'h33f4: o_data_a = 16'b1110110000010000;
            14'h33f5: o_data_a = 16'b0000000000001110;
            14'h33f6: o_data_a = 16'b1110001100001000;
            14'h33f7: o_data_a = 16'b0011001111111011;
            14'h33f8: o_data_a = 16'b1110110000010000;
            14'h33f9: o_data_a = 16'b0000000001011111;
            14'h33fa: o_data_a = 16'b1110101010000111;
            14'h33fb: o_data_a = 16'b0000000000000000;
            14'h33fc: o_data_a = 16'b1111110010101000;
            14'h33fd: o_data_a = 16'b1111110000010000;
            14'h33fe: o_data_a = 16'b0000000000000101;
            14'h33ff: o_data_a = 16'b1110001100001000;
            14'h3400: o_data_a = 16'b0000000001001000;
            14'h3401: o_data_a = 16'b1110110000010000;
            14'h3402: o_data_a = 16'b0000000000000000;
            14'h3403: o_data_a = 16'b1111110111101000;
            14'h3404: o_data_a = 16'b1110110010100000;
            14'h3405: o_data_a = 16'b1110001100001000;
            14'h3406: o_data_a = 16'b0000000000110011;
            14'h3407: o_data_a = 16'b1110110000010000;
            14'h3408: o_data_a = 16'b0000000000000000;
            14'h3409: o_data_a = 16'b1111110111101000;
            14'h340a: o_data_a = 16'b1110110010100000;
            14'h340b: o_data_a = 16'b1110001100001000;
            14'h340c: o_data_a = 16'b0000000000110011;
            14'h340d: o_data_a = 16'b1110110000010000;
            14'h340e: o_data_a = 16'b0000000000000000;
            14'h340f: o_data_a = 16'b1111110111101000;
            14'h3410: o_data_a = 16'b1110110010100000;
            14'h3411: o_data_a = 16'b1110001100001000;
            14'h3412: o_data_a = 16'b0000000000110011;
            14'h3413: o_data_a = 16'b1110110000010000;
            14'h3414: o_data_a = 16'b0000000000000000;
            14'h3415: o_data_a = 16'b1111110111101000;
            14'h3416: o_data_a = 16'b1110110010100000;
            14'h3417: o_data_a = 16'b1110001100001000;
            14'h3418: o_data_a = 16'b0000000000110011;
            14'h3419: o_data_a = 16'b1110110000010000;
            14'h341a: o_data_a = 16'b0000000000000000;
            14'h341b: o_data_a = 16'b1111110111101000;
            14'h341c: o_data_a = 16'b1110110010100000;
            14'h341d: o_data_a = 16'b1110001100001000;
            14'h341e: o_data_a = 16'b0000000000111111;
            14'h341f: o_data_a = 16'b1110110000010000;
            14'h3420: o_data_a = 16'b0000000000000000;
            14'h3421: o_data_a = 16'b1111110111101000;
            14'h3422: o_data_a = 16'b1110110010100000;
            14'h3423: o_data_a = 16'b1110001100001000;
            14'h3424: o_data_a = 16'b0000000000110011;
            14'h3425: o_data_a = 16'b1110110000010000;
            14'h3426: o_data_a = 16'b0000000000000000;
            14'h3427: o_data_a = 16'b1111110111101000;
            14'h3428: o_data_a = 16'b1110110010100000;
            14'h3429: o_data_a = 16'b1110001100001000;
            14'h342a: o_data_a = 16'b0000000000110011;
            14'h342b: o_data_a = 16'b1110110000010000;
            14'h342c: o_data_a = 16'b0000000000000000;
            14'h342d: o_data_a = 16'b1111110111101000;
            14'h342e: o_data_a = 16'b1110110010100000;
            14'h342f: o_data_a = 16'b1110001100001000;
            14'h3430: o_data_a = 16'b0000000000110011;
            14'h3431: o_data_a = 16'b1110110000010000;
            14'h3432: o_data_a = 16'b0000000000000000;
            14'h3433: o_data_a = 16'b1111110111101000;
            14'h3434: o_data_a = 16'b1110110010100000;
            14'h3435: o_data_a = 16'b1110001100001000;
            14'h3436: o_data_a = 16'b0000000000110011;
            14'h3437: o_data_a = 16'b1110110000010000;
            14'h3438: o_data_a = 16'b0000000000000000;
            14'h3439: o_data_a = 16'b1111110111101000;
            14'h343a: o_data_a = 16'b1110110010100000;
            14'h343b: o_data_a = 16'b1110001100001000;
            14'h343c: o_data_a = 16'b0000000000000000;
            14'h343d: o_data_a = 16'b1111110111001000;
            14'h343e: o_data_a = 16'b1111110010100000;
            14'h343f: o_data_a = 16'b1110101010001000;
            14'h3440: o_data_a = 16'b0000000000000000;
            14'h3441: o_data_a = 16'b1111110111001000;
            14'h3442: o_data_a = 16'b1111110010100000;
            14'h3443: o_data_a = 16'b1110101010001000;
            14'h3444: o_data_a = 16'b0000000000001100;
            14'h3445: o_data_a = 16'b1110110000010000;
            14'h3446: o_data_a = 16'b0000000000001101;
            14'h3447: o_data_a = 16'b1110001100001000;
            14'h3448: o_data_a = 16'b0100010110110011;
            14'h3449: o_data_a = 16'b1110110000010000;
            14'h344a: o_data_a = 16'b0000000000001110;
            14'h344b: o_data_a = 16'b1110001100001000;
            14'h344c: o_data_a = 16'b0011010001010000;
            14'h344d: o_data_a = 16'b1110110000010000;
            14'h344e: o_data_a = 16'b0000000001011111;
            14'h344f: o_data_a = 16'b1110101010000111;
            14'h3450: o_data_a = 16'b0000000000000000;
            14'h3451: o_data_a = 16'b1111110010101000;
            14'h3452: o_data_a = 16'b1111110000010000;
            14'h3453: o_data_a = 16'b0000000000000101;
            14'h3454: o_data_a = 16'b1110001100001000;
            14'h3455: o_data_a = 16'b0000000001001001;
            14'h3456: o_data_a = 16'b1110110000010000;
            14'h3457: o_data_a = 16'b0000000000000000;
            14'h3458: o_data_a = 16'b1111110111101000;
            14'h3459: o_data_a = 16'b1110110010100000;
            14'h345a: o_data_a = 16'b1110001100001000;
            14'h345b: o_data_a = 16'b0000000000011110;
            14'h345c: o_data_a = 16'b1110110000010000;
            14'h345d: o_data_a = 16'b0000000000000000;
            14'h345e: o_data_a = 16'b1111110111101000;
            14'h345f: o_data_a = 16'b1110110010100000;
            14'h3460: o_data_a = 16'b1110001100001000;
            14'h3461: o_data_a = 16'b0000000000001100;
            14'h3462: o_data_a = 16'b1110110000010000;
            14'h3463: o_data_a = 16'b0000000000000000;
            14'h3464: o_data_a = 16'b1111110111101000;
            14'h3465: o_data_a = 16'b1110110010100000;
            14'h3466: o_data_a = 16'b1110001100001000;
            14'h3467: o_data_a = 16'b0000000000001100;
            14'h3468: o_data_a = 16'b1110110000010000;
            14'h3469: o_data_a = 16'b0000000000000000;
            14'h346a: o_data_a = 16'b1111110111101000;
            14'h346b: o_data_a = 16'b1110110010100000;
            14'h346c: o_data_a = 16'b1110001100001000;
            14'h346d: o_data_a = 16'b0000000000001100;
            14'h346e: o_data_a = 16'b1110110000010000;
            14'h346f: o_data_a = 16'b0000000000000000;
            14'h3470: o_data_a = 16'b1111110111101000;
            14'h3471: o_data_a = 16'b1110110010100000;
            14'h3472: o_data_a = 16'b1110001100001000;
            14'h3473: o_data_a = 16'b0000000000001100;
            14'h3474: o_data_a = 16'b1110110000010000;
            14'h3475: o_data_a = 16'b0000000000000000;
            14'h3476: o_data_a = 16'b1111110111101000;
            14'h3477: o_data_a = 16'b1110110010100000;
            14'h3478: o_data_a = 16'b1110001100001000;
            14'h3479: o_data_a = 16'b0000000000001100;
            14'h347a: o_data_a = 16'b1110110000010000;
            14'h347b: o_data_a = 16'b0000000000000000;
            14'h347c: o_data_a = 16'b1111110111101000;
            14'h347d: o_data_a = 16'b1110110010100000;
            14'h347e: o_data_a = 16'b1110001100001000;
            14'h347f: o_data_a = 16'b0000000000001100;
            14'h3480: o_data_a = 16'b1110110000010000;
            14'h3481: o_data_a = 16'b0000000000000000;
            14'h3482: o_data_a = 16'b1111110111101000;
            14'h3483: o_data_a = 16'b1110110010100000;
            14'h3484: o_data_a = 16'b1110001100001000;
            14'h3485: o_data_a = 16'b0000000000001100;
            14'h3486: o_data_a = 16'b1110110000010000;
            14'h3487: o_data_a = 16'b0000000000000000;
            14'h3488: o_data_a = 16'b1111110111101000;
            14'h3489: o_data_a = 16'b1110110010100000;
            14'h348a: o_data_a = 16'b1110001100001000;
            14'h348b: o_data_a = 16'b0000000000011110;
            14'h348c: o_data_a = 16'b1110110000010000;
            14'h348d: o_data_a = 16'b0000000000000000;
            14'h348e: o_data_a = 16'b1111110111101000;
            14'h348f: o_data_a = 16'b1110110010100000;
            14'h3490: o_data_a = 16'b1110001100001000;
            14'h3491: o_data_a = 16'b0000000000000000;
            14'h3492: o_data_a = 16'b1111110111001000;
            14'h3493: o_data_a = 16'b1111110010100000;
            14'h3494: o_data_a = 16'b1110101010001000;
            14'h3495: o_data_a = 16'b0000000000000000;
            14'h3496: o_data_a = 16'b1111110111001000;
            14'h3497: o_data_a = 16'b1111110010100000;
            14'h3498: o_data_a = 16'b1110101010001000;
            14'h3499: o_data_a = 16'b0000000000001100;
            14'h349a: o_data_a = 16'b1110110000010000;
            14'h349b: o_data_a = 16'b0000000000001101;
            14'h349c: o_data_a = 16'b1110001100001000;
            14'h349d: o_data_a = 16'b0100010110110011;
            14'h349e: o_data_a = 16'b1110110000010000;
            14'h349f: o_data_a = 16'b0000000000001110;
            14'h34a0: o_data_a = 16'b1110001100001000;
            14'h34a1: o_data_a = 16'b0011010010100101;
            14'h34a2: o_data_a = 16'b1110110000010000;
            14'h34a3: o_data_a = 16'b0000000001011111;
            14'h34a4: o_data_a = 16'b1110101010000111;
            14'h34a5: o_data_a = 16'b0000000000000000;
            14'h34a6: o_data_a = 16'b1111110010101000;
            14'h34a7: o_data_a = 16'b1111110000010000;
            14'h34a8: o_data_a = 16'b0000000000000101;
            14'h34a9: o_data_a = 16'b1110001100001000;
            14'h34aa: o_data_a = 16'b0000000001001010;
            14'h34ab: o_data_a = 16'b1110110000010000;
            14'h34ac: o_data_a = 16'b0000000000000000;
            14'h34ad: o_data_a = 16'b1111110111101000;
            14'h34ae: o_data_a = 16'b1110110010100000;
            14'h34af: o_data_a = 16'b1110001100001000;
            14'h34b0: o_data_a = 16'b0000000000111100;
            14'h34b1: o_data_a = 16'b1110110000010000;
            14'h34b2: o_data_a = 16'b0000000000000000;
            14'h34b3: o_data_a = 16'b1111110111101000;
            14'h34b4: o_data_a = 16'b1110110010100000;
            14'h34b5: o_data_a = 16'b1110001100001000;
            14'h34b6: o_data_a = 16'b0000000000011000;
            14'h34b7: o_data_a = 16'b1110110000010000;
            14'h34b8: o_data_a = 16'b0000000000000000;
            14'h34b9: o_data_a = 16'b1111110111101000;
            14'h34ba: o_data_a = 16'b1110110010100000;
            14'h34bb: o_data_a = 16'b1110001100001000;
            14'h34bc: o_data_a = 16'b0000000000011000;
            14'h34bd: o_data_a = 16'b1110110000010000;
            14'h34be: o_data_a = 16'b0000000000000000;
            14'h34bf: o_data_a = 16'b1111110111101000;
            14'h34c0: o_data_a = 16'b1110110010100000;
            14'h34c1: o_data_a = 16'b1110001100001000;
            14'h34c2: o_data_a = 16'b0000000000011000;
            14'h34c3: o_data_a = 16'b1110110000010000;
            14'h34c4: o_data_a = 16'b0000000000000000;
            14'h34c5: o_data_a = 16'b1111110111101000;
            14'h34c6: o_data_a = 16'b1110110010100000;
            14'h34c7: o_data_a = 16'b1110001100001000;
            14'h34c8: o_data_a = 16'b0000000000011000;
            14'h34c9: o_data_a = 16'b1110110000010000;
            14'h34ca: o_data_a = 16'b0000000000000000;
            14'h34cb: o_data_a = 16'b1111110111101000;
            14'h34cc: o_data_a = 16'b1110110010100000;
            14'h34cd: o_data_a = 16'b1110001100001000;
            14'h34ce: o_data_a = 16'b0000000000011000;
            14'h34cf: o_data_a = 16'b1110110000010000;
            14'h34d0: o_data_a = 16'b0000000000000000;
            14'h34d1: o_data_a = 16'b1111110111101000;
            14'h34d2: o_data_a = 16'b1110110010100000;
            14'h34d3: o_data_a = 16'b1110001100001000;
            14'h34d4: o_data_a = 16'b0000000000011011;
            14'h34d5: o_data_a = 16'b1110110000010000;
            14'h34d6: o_data_a = 16'b0000000000000000;
            14'h34d7: o_data_a = 16'b1111110111101000;
            14'h34d8: o_data_a = 16'b1110110010100000;
            14'h34d9: o_data_a = 16'b1110001100001000;
            14'h34da: o_data_a = 16'b0000000000011011;
            14'h34db: o_data_a = 16'b1110110000010000;
            14'h34dc: o_data_a = 16'b0000000000000000;
            14'h34dd: o_data_a = 16'b1111110111101000;
            14'h34de: o_data_a = 16'b1110110010100000;
            14'h34df: o_data_a = 16'b1110001100001000;
            14'h34e0: o_data_a = 16'b0000000000001110;
            14'h34e1: o_data_a = 16'b1110110000010000;
            14'h34e2: o_data_a = 16'b0000000000000000;
            14'h34e3: o_data_a = 16'b1111110111101000;
            14'h34e4: o_data_a = 16'b1110110010100000;
            14'h34e5: o_data_a = 16'b1110001100001000;
            14'h34e6: o_data_a = 16'b0000000000000000;
            14'h34e7: o_data_a = 16'b1111110111001000;
            14'h34e8: o_data_a = 16'b1111110010100000;
            14'h34e9: o_data_a = 16'b1110101010001000;
            14'h34ea: o_data_a = 16'b0000000000000000;
            14'h34eb: o_data_a = 16'b1111110111001000;
            14'h34ec: o_data_a = 16'b1111110010100000;
            14'h34ed: o_data_a = 16'b1110101010001000;
            14'h34ee: o_data_a = 16'b0000000000001100;
            14'h34ef: o_data_a = 16'b1110110000010000;
            14'h34f0: o_data_a = 16'b0000000000001101;
            14'h34f1: o_data_a = 16'b1110001100001000;
            14'h34f2: o_data_a = 16'b0100010110110011;
            14'h34f3: o_data_a = 16'b1110110000010000;
            14'h34f4: o_data_a = 16'b0000000000001110;
            14'h34f5: o_data_a = 16'b1110001100001000;
            14'h34f6: o_data_a = 16'b0011010011111010;
            14'h34f7: o_data_a = 16'b1110110000010000;
            14'h34f8: o_data_a = 16'b0000000001011111;
            14'h34f9: o_data_a = 16'b1110101010000111;
            14'h34fa: o_data_a = 16'b0000000000000000;
            14'h34fb: o_data_a = 16'b1111110010101000;
            14'h34fc: o_data_a = 16'b1111110000010000;
            14'h34fd: o_data_a = 16'b0000000000000101;
            14'h34fe: o_data_a = 16'b1110001100001000;
            14'h34ff: o_data_a = 16'b0000000001001011;
            14'h3500: o_data_a = 16'b1110110000010000;
            14'h3501: o_data_a = 16'b0000000000000000;
            14'h3502: o_data_a = 16'b1111110111101000;
            14'h3503: o_data_a = 16'b1110110010100000;
            14'h3504: o_data_a = 16'b1110001100001000;
            14'h3505: o_data_a = 16'b0000000000110011;
            14'h3506: o_data_a = 16'b1110110000010000;
            14'h3507: o_data_a = 16'b0000000000000000;
            14'h3508: o_data_a = 16'b1111110111101000;
            14'h3509: o_data_a = 16'b1110110010100000;
            14'h350a: o_data_a = 16'b1110001100001000;
            14'h350b: o_data_a = 16'b0000000000110011;
            14'h350c: o_data_a = 16'b1110110000010000;
            14'h350d: o_data_a = 16'b0000000000000000;
            14'h350e: o_data_a = 16'b1111110111101000;
            14'h350f: o_data_a = 16'b1110110010100000;
            14'h3510: o_data_a = 16'b1110001100001000;
            14'h3511: o_data_a = 16'b0000000000110011;
            14'h3512: o_data_a = 16'b1110110000010000;
            14'h3513: o_data_a = 16'b0000000000000000;
            14'h3514: o_data_a = 16'b1111110111101000;
            14'h3515: o_data_a = 16'b1110110010100000;
            14'h3516: o_data_a = 16'b1110001100001000;
            14'h3517: o_data_a = 16'b0000000000011011;
            14'h3518: o_data_a = 16'b1110110000010000;
            14'h3519: o_data_a = 16'b0000000000000000;
            14'h351a: o_data_a = 16'b1111110111101000;
            14'h351b: o_data_a = 16'b1110110010100000;
            14'h351c: o_data_a = 16'b1110001100001000;
            14'h351d: o_data_a = 16'b0000000000001111;
            14'h351e: o_data_a = 16'b1110110000010000;
            14'h351f: o_data_a = 16'b0000000000000000;
            14'h3520: o_data_a = 16'b1111110111101000;
            14'h3521: o_data_a = 16'b1110110010100000;
            14'h3522: o_data_a = 16'b1110001100001000;
            14'h3523: o_data_a = 16'b0000000000011011;
            14'h3524: o_data_a = 16'b1110110000010000;
            14'h3525: o_data_a = 16'b0000000000000000;
            14'h3526: o_data_a = 16'b1111110111101000;
            14'h3527: o_data_a = 16'b1110110010100000;
            14'h3528: o_data_a = 16'b1110001100001000;
            14'h3529: o_data_a = 16'b0000000000110011;
            14'h352a: o_data_a = 16'b1110110000010000;
            14'h352b: o_data_a = 16'b0000000000000000;
            14'h352c: o_data_a = 16'b1111110111101000;
            14'h352d: o_data_a = 16'b1110110010100000;
            14'h352e: o_data_a = 16'b1110001100001000;
            14'h352f: o_data_a = 16'b0000000000110011;
            14'h3530: o_data_a = 16'b1110110000010000;
            14'h3531: o_data_a = 16'b0000000000000000;
            14'h3532: o_data_a = 16'b1111110111101000;
            14'h3533: o_data_a = 16'b1110110010100000;
            14'h3534: o_data_a = 16'b1110001100001000;
            14'h3535: o_data_a = 16'b0000000000110011;
            14'h3536: o_data_a = 16'b1110110000010000;
            14'h3537: o_data_a = 16'b0000000000000000;
            14'h3538: o_data_a = 16'b1111110111101000;
            14'h3539: o_data_a = 16'b1110110010100000;
            14'h353a: o_data_a = 16'b1110001100001000;
            14'h353b: o_data_a = 16'b0000000000000000;
            14'h353c: o_data_a = 16'b1111110111001000;
            14'h353d: o_data_a = 16'b1111110010100000;
            14'h353e: o_data_a = 16'b1110101010001000;
            14'h353f: o_data_a = 16'b0000000000000000;
            14'h3540: o_data_a = 16'b1111110111001000;
            14'h3541: o_data_a = 16'b1111110010100000;
            14'h3542: o_data_a = 16'b1110101010001000;
            14'h3543: o_data_a = 16'b0000000000001100;
            14'h3544: o_data_a = 16'b1110110000010000;
            14'h3545: o_data_a = 16'b0000000000001101;
            14'h3546: o_data_a = 16'b1110001100001000;
            14'h3547: o_data_a = 16'b0100010110110011;
            14'h3548: o_data_a = 16'b1110110000010000;
            14'h3549: o_data_a = 16'b0000000000001110;
            14'h354a: o_data_a = 16'b1110001100001000;
            14'h354b: o_data_a = 16'b0011010101001111;
            14'h354c: o_data_a = 16'b1110110000010000;
            14'h354d: o_data_a = 16'b0000000001011111;
            14'h354e: o_data_a = 16'b1110101010000111;
            14'h354f: o_data_a = 16'b0000000000000000;
            14'h3550: o_data_a = 16'b1111110010101000;
            14'h3551: o_data_a = 16'b1111110000010000;
            14'h3552: o_data_a = 16'b0000000000000101;
            14'h3553: o_data_a = 16'b1110001100001000;
            14'h3554: o_data_a = 16'b0000000001001100;
            14'h3555: o_data_a = 16'b1110110000010000;
            14'h3556: o_data_a = 16'b0000000000000000;
            14'h3557: o_data_a = 16'b1111110111101000;
            14'h3558: o_data_a = 16'b1110110010100000;
            14'h3559: o_data_a = 16'b1110001100001000;
            14'h355a: o_data_a = 16'b0000000000000011;
            14'h355b: o_data_a = 16'b1110110000010000;
            14'h355c: o_data_a = 16'b0000000000000000;
            14'h355d: o_data_a = 16'b1111110111101000;
            14'h355e: o_data_a = 16'b1110110010100000;
            14'h355f: o_data_a = 16'b1110001100001000;
            14'h3560: o_data_a = 16'b0000000000000011;
            14'h3561: o_data_a = 16'b1110110000010000;
            14'h3562: o_data_a = 16'b0000000000000000;
            14'h3563: o_data_a = 16'b1111110111101000;
            14'h3564: o_data_a = 16'b1110110010100000;
            14'h3565: o_data_a = 16'b1110001100001000;
            14'h3566: o_data_a = 16'b0000000000000011;
            14'h3567: o_data_a = 16'b1110110000010000;
            14'h3568: o_data_a = 16'b0000000000000000;
            14'h3569: o_data_a = 16'b1111110111101000;
            14'h356a: o_data_a = 16'b1110110010100000;
            14'h356b: o_data_a = 16'b1110001100001000;
            14'h356c: o_data_a = 16'b0000000000000011;
            14'h356d: o_data_a = 16'b1110110000010000;
            14'h356e: o_data_a = 16'b0000000000000000;
            14'h356f: o_data_a = 16'b1111110111101000;
            14'h3570: o_data_a = 16'b1110110010100000;
            14'h3571: o_data_a = 16'b1110001100001000;
            14'h3572: o_data_a = 16'b0000000000000011;
            14'h3573: o_data_a = 16'b1110110000010000;
            14'h3574: o_data_a = 16'b0000000000000000;
            14'h3575: o_data_a = 16'b1111110111101000;
            14'h3576: o_data_a = 16'b1110110010100000;
            14'h3577: o_data_a = 16'b1110001100001000;
            14'h3578: o_data_a = 16'b0000000000000011;
            14'h3579: o_data_a = 16'b1110110000010000;
            14'h357a: o_data_a = 16'b0000000000000000;
            14'h357b: o_data_a = 16'b1111110111101000;
            14'h357c: o_data_a = 16'b1110110010100000;
            14'h357d: o_data_a = 16'b1110001100001000;
            14'h357e: o_data_a = 16'b0000000000100011;
            14'h357f: o_data_a = 16'b1110110000010000;
            14'h3580: o_data_a = 16'b0000000000000000;
            14'h3581: o_data_a = 16'b1111110111101000;
            14'h3582: o_data_a = 16'b1110110010100000;
            14'h3583: o_data_a = 16'b1110001100001000;
            14'h3584: o_data_a = 16'b0000000000110011;
            14'h3585: o_data_a = 16'b1110110000010000;
            14'h3586: o_data_a = 16'b0000000000000000;
            14'h3587: o_data_a = 16'b1111110111101000;
            14'h3588: o_data_a = 16'b1110110010100000;
            14'h3589: o_data_a = 16'b1110001100001000;
            14'h358a: o_data_a = 16'b0000000000111111;
            14'h358b: o_data_a = 16'b1110110000010000;
            14'h358c: o_data_a = 16'b0000000000000000;
            14'h358d: o_data_a = 16'b1111110111101000;
            14'h358e: o_data_a = 16'b1110110010100000;
            14'h358f: o_data_a = 16'b1110001100001000;
            14'h3590: o_data_a = 16'b0000000000000000;
            14'h3591: o_data_a = 16'b1111110111001000;
            14'h3592: o_data_a = 16'b1111110010100000;
            14'h3593: o_data_a = 16'b1110101010001000;
            14'h3594: o_data_a = 16'b0000000000000000;
            14'h3595: o_data_a = 16'b1111110111001000;
            14'h3596: o_data_a = 16'b1111110010100000;
            14'h3597: o_data_a = 16'b1110101010001000;
            14'h3598: o_data_a = 16'b0000000000001100;
            14'h3599: o_data_a = 16'b1110110000010000;
            14'h359a: o_data_a = 16'b0000000000001101;
            14'h359b: o_data_a = 16'b1110001100001000;
            14'h359c: o_data_a = 16'b0100010110110011;
            14'h359d: o_data_a = 16'b1110110000010000;
            14'h359e: o_data_a = 16'b0000000000001110;
            14'h359f: o_data_a = 16'b1110001100001000;
            14'h35a0: o_data_a = 16'b0011010110100100;
            14'h35a1: o_data_a = 16'b1110110000010000;
            14'h35a2: o_data_a = 16'b0000000001011111;
            14'h35a3: o_data_a = 16'b1110101010000111;
            14'h35a4: o_data_a = 16'b0000000000000000;
            14'h35a5: o_data_a = 16'b1111110010101000;
            14'h35a6: o_data_a = 16'b1111110000010000;
            14'h35a7: o_data_a = 16'b0000000000000101;
            14'h35a8: o_data_a = 16'b1110001100001000;
            14'h35a9: o_data_a = 16'b0000000001001101;
            14'h35aa: o_data_a = 16'b1110110000010000;
            14'h35ab: o_data_a = 16'b0000000000000000;
            14'h35ac: o_data_a = 16'b1111110111101000;
            14'h35ad: o_data_a = 16'b1110110010100000;
            14'h35ae: o_data_a = 16'b1110001100001000;
            14'h35af: o_data_a = 16'b0000000000100001;
            14'h35b0: o_data_a = 16'b1110110000010000;
            14'h35b1: o_data_a = 16'b0000000000000000;
            14'h35b2: o_data_a = 16'b1111110111101000;
            14'h35b3: o_data_a = 16'b1110110010100000;
            14'h35b4: o_data_a = 16'b1110001100001000;
            14'h35b5: o_data_a = 16'b0000000000110011;
            14'h35b6: o_data_a = 16'b1110110000010000;
            14'h35b7: o_data_a = 16'b0000000000000000;
            14'h35b8: o_data_a = 16'b1111110111101000;
            14'h35b9: o_data_a = 16'b1110110010100000;
            14'h35ba: o_data_a = 16'b1110001100001000;
            14'h35bb: o_data_a = 16'b0000000000111111;
            14'h35bc: o_data_a = 16'b1110110000010000;
            14'h35bd: o_data_a = 16'b0000000000000000;
            14'h35be: o_data_a = 16'b1111110111101000;
            14'h35bf: o_data_a = 16'b1110110010100000;
            14'h35c0: o_data_a = 16'b1110001100001000;
            14'h35c1: o_data_a = 16'b0000000000111111;
            14'h35c2: o_data_a = 16'b1110110000010000;
            14'h35c3: o_data_a = 16'b0000000000000000;
            14'h35c4: o_data_a = 16'b1111110111101000;
            14'h35c5: o_data_a = 16'b1110110010100000;
            14'h35c6: o_data_a = 16'b1110001100001000;
            14'h35c7: o_data_a = 16'b0000000000110011;
            14'h35c8: o_data_a = 16'b1110110000010000;
            14'h35c9: o_data_a = 16'b0000000000000000;
            14'h35ca: o_data_a = 16'b1111110111101000;
            14'h35cb: o_data_a = 16'b1110110010100000;
            14'h35cc: o_data_a = 16'b1110001100001000;
            14'h35cd: o_data_a = 16'b0000000000110011;
            14'h35ce: o_data_a = 16'b1110110000010000;
            14'h35cf: o_data_a = 16'b0000000000000000;
            14'h35d0: o_data_a = 16'b1111110111101000;
            14'h35d1: o_data_a = 16'b1110110010100000;
            14'h35d2: o_data_a = 16'b1110001100001000;
            14'h35d3: o_data_a = 16'b0000000000110011;
            14'h35d4: o_data_a = 16'b1110110000010000;
            14'h35d5: o_data_a = 16'b0000000000000000;
            14'h35d6: o_data_a = 16'b1111110111101000;
            14'h35d7: o_data_a = 16'b1110110010100000;
            14'h35d8: o_data_a = 16'b1110001100001000;
            14'h35d9: o_data_a = 16'b0000000000110011;
            14'h35da: o_data_a = 16'b1110110000010000;
            14'h35db: o_data_a = 16'b0000000000000000;
            14'h35dc: o_data_a = 16'b1111110111101000;
            14'h35dd: o_data_a = 16'b1110110010100000;
            14'h35de: o_data_a = 16'b1110001100001000;
            14'h35df: o_data_a = 16'b0000000000110011;
            14'h35e0: o_data_a = 16'b1110110000010000;
            14'h35e1: o_data_a = 16'b0000000000000000;
            14'h35e2: o_data_a = 16'b1111110111101000;
            14'h35e3: o_data_a = 16'b1110110010100000;
            14'h35e4: o_data_a = 16'b1110001100001000;
            14'h35e5: o_data_a = 16'b0000000000000000;
            14'h35e6: o_data_a = 16'b1111110111001000;
            14'h35e7: o_data_a = 16'b1111110010100000;
            14'h35e8: o_data_a = 16'b1110101010001000;
            14'h35e9: o_data_a = 16'b0000000000000000;
            14'h35ea: o_data_a = 16'b1111110111001000;
            14'h35eb: o_data_a = 16'b1111110010100000;
            14'h35ec: o_data_a = 16'b1110101010001000;
            14'h35ed: o_data_a = 16'b0000000000001100;
            14'h35ee: o_data_a = 16'b1110110000010000;
            14'h35ef: o_data_a = 16'b0000000000001101;
            14'h35f0: o_data_a = 16'b1110001100001000;
            14'h35f1: o_data_a = 16'b0100010110110011;
            14'h35f2: o_data_a = 16'b1110110000010000;
            14'h35f3: o_data_a = 16'b0000000000001110;
            14'h35f4: o_data_a = 16'b1110001100001000;
            14'h35f5: o_data_a = 16'b0011010111111001;
            14'h35f6: o_data_a = 16'b1110110000010000;
            14'h35f7: o_data_a = 16'b0000000001011111;
            14'h35f8: o_data_a = 16'b1110101010000111;
            14'h35f9: o_data_a = 16'b0000000000000000;
            14'h35fa: o_data_a = 16'b1111110010101000;
            14'h35fb: o_data_a = 16'b1111110000010000;
            14'h35fc: o_data_a = 16'b0000000000000101;
            14'h35fd: o_data_a = 16'b1110001100001000;
            14'h35fe: o_data_a = 16'b0000000001001110;
            14'h35ff: o_data_a = 16'b1110110000010000;
            14'h3600: o_data_a = 16'b0000000000000000;
            14'h3601: o_data_a = 16'b1111110111101000;
            14'h3602: o_data_a = 16'b1110110010100000;
            14'h3603: o_data_a = 16'b1110001100001000;
            14'h3604: o_data_a = 16'b0000000000110011;
            14'h3605: o_data_a = 16'b1110110000010000;
            14'h3606: o_data_a = 16'b0000000000000000;
            14'h3607: o_data_a = 16'b1111110111101000;
            14'h3608: o_data_a = 16'b1110110010100000;
            14'h3609: o_data_a = 16'b1110001100001000;
            14'h360a: o_data_a = 16'b0000000000110011;
            14'h360b: o_data_a = 16'b1110110000010000;
            14'h360c: o_data_a = 16'b0000000000000000;
            14'h360d: o_data_a = 16'b1111110111101000;
            14'h360e: o_data_a = 16'b1110110010100000;
            14'h360f: o_data_a = 16'b1110001100001000;
            14'h3610: o_data_a = 16'b0000000000110111;
            14'h3611: o_data_a = 16'b1110110000010000;
            14'h3612: o_data_a = 16'b0000000000000000;
            14'h3613: o_data_a = 16'b1111110111101000;
            14'h3614: o_data_a = 16'b1110110010100000;
            14'h3615: o_data_a = 16'b1110001100001000;
            14'h3616: o_data_a = 16'b0000000000110111;
            14'h3617: o_data_a = 16'b1110110000010000;
            14'h3618: o_data_a = 16'b0000000000000000;
            14'h3619: o_data_a = 16'b1111110111101000;
            14'h361a: o_data_a = 16'b1110110010100000;
            14'h361b: o_data_a = 16'b1110001100001000;
            14'h361c: o_data_a = 16'b0000000000111111;
            14'h361d: o_data_a = 16'b1110110000010000;
            14'h361e: o_data_a = 16'b0000000000000000;
            14'h361f: o_data_a = 16'b1111110111101000;
            14'h3620: o_data_a = 16'b1110110010100000;
            14'h3621: o_data_a = 16'b1110001100001000;
            14'h3622: o_data_a = 16'b0000000000111011;
            14'h3623: o_data_a = 16'b1110110000010000;
            14'h3624: o_data_a = 16'b0000000000000000;
            14'h3625: o_data_a = 16'b1111110111101000;
            14'h3626: o_data_a = 16'b1110110010100000;
            14'h3627: o_data_a = 16'b1110001100001000;
            14'h3628: o_data_a = 16'b0000000000111011;
            14'h3629: o_data_a = 16'b1110110000010000;
            14'h362a: o_data_a = 16'b0000000000000000;
            14'h362b: o_data_a = 16'b1111110111101000;
            14'h362c: o_data_a = 16'b1110110010100000;
            14'h362d: o_data_a = 16'b1110001100001000;
            14'h362e: o_data_a = 16'b0000000000110011;
            14'h362f: o_data_a = 16'b1110110000010000;
            14'h3630: o_data_a = 16'b0000000000000000;
            14'h3631: o_data_a = 16'b1111110111101000;
            14'h3632: o_data_a = 16'b1110110010100000;
            14'h3633: o_data_a = 16'b1110001100001000;
            14'h3634: o_data_a = 16'b0000000000110011;
            14'h3635: o_data_a = 16'b1110110000010000;
            14'h3636: o_data_a = 16'b0000000000000000;
            14'h3637: o_data_a = 16'b1111110111101000;
            14'h3638: o_data_a = 16'b1110110010100000;
            14'h3639: o_data_a = 16'b1110001100001000;
            14'h363a: o_data_a = 16'b0000000000000000;
            14'h363b: o_data_a = 16'b1111110111001000;
            14'h363c: o_data_a = 16'b1111110010100000;
            14'h363d: o_data_a = 16'b1110101010001000;
            14'h363e: o_data_a = 16'b0000000000000000;
            14'h363f: o_data_a = 16'b1111110111001000;
            14'h3640: o_data_a = 16'b1111110010100000;
            14'h3641: o_data_a = 16'b1110101010001000;
            14'h3642: o_data_a = 16'b0000000000001100;
            14'h3643: o_data_a = 16'b1110110000010000;
            14'h3644: o_data_a = 16'b0000000000001101;
            14'h3645: o_data_a = 16'b1110001100001000;
            14'h3646: o_data_a = 16'b0100010110110011;
            14'h3647: o_data_a = 16'b1110110000010000;
            14'h3648: o_data_a = 16'b0000000000001110;
            14'h3649: o_data_a = 16'b1110001100001000;
            14'h364a: o_data_a = 16'b0011011001001110;
            14'h364b: o_data_a = 16'b1110110000010000;
            14'h364c: o_data_a = 16'b0000000001011111;
            14'h364d: o_data_a = 16'b1110101010000111;
            14'h364e: o_data_a = 16'b0000000000000000;
            14'h364f: o_data_a = 16'b1111110010101000;
            14'h3650: o_data_a = 16'b1111110000010000;
            14'h3651: o_data_a = 16'b0000000000000101;
            14'h3652: o_data_a = 16'b1110001100001000;
            14'h3653: o_data_a = 16'b0000000001001111;
            14'h3654: o_data_a = 16'b1110110000010000;
            14'h3655: o_data_a = 16'b0000000000000000;
            14'h3656: o_data_a = 16'b1111110111101000;
            14'h3657: o_data_a = 16'b1110110010100000;
            14'h3658: o_data_a = 16'b1110001100001000;
            14'h3659: o_data_a = 16'b0000000000011110;
            14'h365a: o_data_a = 16'b1110110000010000;
            14'h365b: o_data_a = 16'b0000000000000000;
            14'h365c: o_data_a = 16'b1111110111101000;
            14'h365d: o_data_a = 16'b1110110010100000;
            14'h365e: o_data_a = 16'b1110001100001000;
            14'h365f: o_data_a = 16'b0000000000110011;
            14'h3660: o_data_a = 16'b1110110000010000;
            14'h3661: o_data_a = 16'b0000000000000000;
            14'h3662: o_data_a = 16'b1111110111101000;
            14'h3663: o_data_a = 16'b1110110010100000;
            14'h3664: o_data_a = 16'b1110001100001000;
            14'h3665: o_data_a = 16'b0000000000110011;
            14'h3666: o_data_a = 16'b1110110000010000;
            14'h3667: o_data_a = 16'b0000000000000000;
            14'h3668: o_data_a = 16'b1111110111101000;
            14'h3669: o_data_a = 16'b1110110010100000;
            14'h366a: o_data_a = 16'b1110001100001000;
            14'h366b: o_data_a = 16'b0000000000110011;
            14'h366c: o_data_a = 16'b1110110000010000;
            14'h366d: o_data_a = 16'b0000000000000000;
            14'h366e: o_data_a = 16'b1111110111101000;
            14'h366f: o_data_a = 16'b1110110010100000;
            14'h3670: o_data_a = 16'b1110001100001000;
            14'h3671: o_data_a = 16'b0000000000110011;
            14'h3672: o_data_a = 16'b1110110000010000;
            14'h3673: o_data_a = 16'b0000000000000000;
            14'h3674: o_data_a = 16'b1111110111101000;
            14'h3675: o_data_a = 16'b1110110010100000;
            14'h3676: o_data_a = 16'b1110001100001000;
            14'h3677: o_data_a = 16'b0000000000110011;
            14'h3678: o_data_a = 16'b1110110000010000;
            14'h3679: o_data_a = 16'b0000000000000000;
            14'h367a: o_data_a = 16'b1111110111101000;
            14'h367b: o_data_a = 16'b1110110010100000;
            14'h367c: o_data_a = 16'b1110001100001000;
            14'h367d: o_data_a = 16'b0000000000110011;
            14'h367e: o_data_a = 16'b1110110000010000;
            14'h367f: o_data_a = 16'b0000000000000000;
            14'h3680: o_data_a = 16'b1111110111101000;
            14'h3681: o_data_a = 16'b1110110010100000;
            14'h3682: o_data_a = 16'b1110001100001000;
            14'h3683: o_data_a = 16'b0000000000110011;
            14'h3684: o_data_a = 16'b1110110000010000;
            14'h3685: o_data_a = 16'b0000000000000000;
            14'h3686: o_data_a = 16'b1111110111101000;
            14'h3687: o_data_a = 16'b1110110010100000;
            14'h3688: o_data_a = 16'b1110001100001000;
            14'h3689: o_data_a = 16'b0000000000011110;
            14'h368a: o_data_a = 16'b1110110000010000;
            14'h368b: o_data_a = 16'b0000000000000000;
            14'h368c: o_data_a = 16'b1111110111101000;
            14'h368d: o_data_a = 16'b1110110010100000;
            14'h368e: o_data_a = 16'b1110001100001000;
            14'h368f: o_data_a = 16'b0000000000000000;
            14'h3690: o_data_a = 16'b1111110111001000;
            14'h3691: o_data_a = 16'b1111110010100000;
            14'h3692: o_data_a = 16'b1110101010001000;
            14'h3693: o_data_a = 16'b0000000000000000;
            14'h3694: o_data_a = 16'b1111110111001000;
            14'h3695: o_data_a = 16'b1111110010100000;
            14'h3696: o_data_a = 16'b1110101010001000;
            14'h3697: o_data_a = 16'b0000000000001100;
            14'h3698: o_data_a = 16'b1110110000010000;
            14'h3699: o_data_a = 16'b0000000000001101;
            14'h369a: o_data_a = 16'b1110001100001000;
            14'h369b: o_data_a = 16'b0100010110110011;
            14'h369c: o_data_a = 16'b1110110000010000;
            14'h369d: o_data_a = 16'b0000000000001110;
            14'h369e: o_data_a = 16'b1110001100001000;
            14'h369f: o_data_a = 16'b0011011010100011;
            14'h36a0: o_data_a = 16'b1110110000010000;
            14'h36a1: o_data_a = 16'b0000000001011111;
            14'h36a2: o_data_a = 16'b1110101010000111;
            14'h36a3: o_data_a = 16'b0000000000000000;
            14'h36a4: o_data_a = 16'b1111110010101000;
            14'h36a5: o_data_a = 16'b1111110000010000;
            14'h36a6: o_data_a = 16'b0000000000000101;
            14'h36a7: o_data_a = 16'b1110001100001000;
            14'h36a8: o_data_a = 16'b0000000001010000;
            14'h36a9: o_data_a = 16'b1110110000010000;
            14'h36aa: o_data_a = 16'b0000000000000000;
            14'h36ab: o_data_a = 16'b1111110111101000;
            14'h36ac: o_data_a = 16'b1110110010100000;
            14'h36ad: o_data_a = 16'b1110001100001000;
            14'h36ae: o_data_a = 16'b0000000000011111;
            14'h36af: o_data_a = 16'b1110110000010000;
            14'h36b0: o_data_a = 16'b0000000000000000;
            14'h36b1: o_data_a = 16'b1111110111101000;
            14'h36b2: o_data_a = 16'b1110110010100000;
            14'h36b3: o_data_a = 16'b1110001100001000;
            14'h36b4: o_data_a = 16'b0000000000110011;
            14'h36b5: o_data_a = 16'b1110110000010000;
            14'h36b6: o_data_a = 16'b0000000000000000;
            14'h36b7: o_data_a = 16'b1111110111101000;
            14'h36b8: o_data_a = 16'b1110110010100000;
            14'h36b9: o_data_a = 16'b1110001100001000;
            14'h36ba: o_data_a = 16'b0000000000110011;
            14'h36bb: o_data_a = 16'b1110110000010000;
            14'h36bc: o_data_a = 16'b0000000000000000;
            14'h36bd: o_data_a = 16'b1111110111101000;
            14'h36be: o_data_a = 16'b1110110010100000;
            14'h36bf: o_data_a = 16'b1110001100001000;
            14'h36c0: o_data_a = 16'b0000000000110011;
            14'h36c1: o_data_a = 16'b1110110000010000;
            14'h36c2: o_data_a = 16'b0000000000000000;
            14'h36c3: o_data_a = 16'b1111110111101000;
            14'h36c4: o_data_a = 16'b1110110010100000;
            14'h36c5: o_data_a = 16'b1110001100001000;
            14'h36c6: o_data_a = 16'b0000000000011111;
            14'h36c7: o_data_a = 16'b1110110000010000;
            14'h36c8: o_data_a = 16'b0000000000000000;
            14'h36c9: o_data_a = 16'b1111110111101000;
            14'h36ca: o_data_a = 16'b1110110010100000;
            14'h36cb: o_data_a = 16'b1110001100001000;
            14'h36cc: o_data_a = 16'b0000000000000011;
            14'h36cd: o_data_a = 16'b1110110000010000;
            14'h36ce: o_data_a = 16'b0000000000000000;
            14'h36cf: o_data_a = 16'b1111110111101000;
            14'h36d0: o_data_a = 16'b1110110010100000;
            14'h36d1: o_data_a = 16'b1110001100001000;
            14'h36d2: o_data_a = 16'b0000000000000011;
            14'h36d3: o_data_a = 16'b1110110000010000;
            14'h36d4: o_data_a = 16'b0000000000000000;
            14'h36d5: o_data_a = 16'b1111110111101000;
            14'h36d6: o_data_a = 16'b1110110010100000;
            14'h36d7: o_data_a = 16'b1110001100001000;
            14'h36d8: o_data_a = 16'b0000000000000011;
            14'h36d9: o_data_a = 16'b1110110000010000;
            14'h36da: o_data_a = 16'b0000000000000000;
            14'h36db: o_data_a = 16'b1111110111101000;
            14'h36dc: o_data_a = 16'b1110110010100000;
            14'h36dd: o_data_a = 16'b1110001100001000;
            14'h36de: o_data_a = 16'b0000000000000011;
            14'h36df: o_data_a = 16'b1110110000010000;
            14'h36e0: o_data_a = 16'b0000000000000000;
            14'h36e1: o_data_a = 16'b1111110111101000;
            14'h36e2: o_data_a = 16'b1110110010100000;
            14'h36e3: o_data_a = 16'b1110001100001000;
            14'h36e4: o_data_a = 16'b0000000000000000;
            14'h36e5: o_data_a = 16'b1111110111001000;
            14'h36e6: o_data_a = 16'b1111110010100000;
            14'h36e7: o_data_a = 16'b1110101010001000;
            14'h36e8: o_data_a = 16'b0000000000000000;
            14'h36e9: o_data_a = 16'b1111110111001000;
            14'h36ea: o_data_a = 16'b1111110010100000;
            14'h36eb: o_data_a = 16'b1110101010001000;
            14'h36ec: o_data_a = 16'b0000000000001100;
            14'h36ed: o_data_a = 16'b1110110000010000;
            14'h36ee: o_data_a = 16'b0000000000001101;
            14'h36ef: o_data_a = 16'b1110001100001000;
            14'h36f0: o_data_a = 16'b0100010110110011;
            14'h36f1: o_data_a = 16'b1110110000010000;
            14'h36f2: o_data_a = 16'b0000000000001110;
            14'h36f3: o_data_a = 16'b1110001100001000;
            14'h36f4: o_data_a = 16'b0011011011111000;
            14'h36f5: o_data_a = 16'b1110110000010000;
            14'h36f6: o_data_a = 16'b0000000001011111;
            14'h36f7: o_data_a = 16'b1110101010000111;
            14'h36f8: o_data_a = 16'b0000000000000000;
            14'h36f9: o_data_a = 16'b1111110010101000;
            14'h36fa: o_data_a = 16'b1111110000010000;
            14'h36fb: o_data_a = 16'b0000000000000101;
            14'h36fc: o_data_a = 16'b1110001100001000;
            14'h36fd: o_data_a = 16'b0000000001010001;
            14'h36fe: o_data_a = 16'b1110110000010000;
            14'h36ff: o_data_a = 16'b0000000000000000;
            14'h3700: o_data_a = 16'b1111110111101000;
            14'h3701: o_data_a = 16'b1110110010100000;
            14'h3702: o_data_a = 16'b1110001100001000;
            14'h3703: o_data_a = 16'b0000000000011110;
            14'h3704: o_data_a = 16'b1110110000010000;
            14'h3705: o_data_a = 16'b0000000000000000;
            14'h3706: o_data_a = 16'b1111110111101000;
            14'h3707: o_data_a = 16'b1110110010100000;
            14'h3708: o_data_a = 16'b1110001100001000;
            14'h3709: o_data_a = 16'b0000000000110011;
            14'h370a: o_data_a = 16'b1110110000010000;
            14'h370b: o_data_a = 16'b0000000000000000;
            14'h370c: o_data_a = 16'b1111110111101000;
            14'h370d: o_data_a = 16'b1110110010100000;
            14'h370e: o_data_a = 16'b1110001100001000;
            14'h370f: o_data_a = 16'b0000000000110011;
            14'h3710: o_data_a = 16'b1110110000010000;
            14'h3711: o_data_a = 16'b0000000000000000;
            14'h3712: o_data_a = 16'b1111110111101000;
            14'h3713: o_data_a = 16'b1110110010100000;
            14'h3714: o_data_a = 16'b1110001100001000;
            14'h3715: o_data_a = 16'b0000000000110011;
            14'h3716: o_data_a = 16'b1110110000010000;
            14'h3717: o_data_a = 16'b0000000000000000;
            14'h3718: o_data_a = 16'b1111110111101000;
            14'h3719: o_data_a = 16'b1110110010100000;
            14'h371a: o_data_a = 16'b1110001100001000;
            14'h371b: o_data_a = 16'b0000000000110011;
            14'h371c: o_data_a = 16'b1110110000010000;
            14'h371d: o_data_a = 16'b0000000000000000;
            14'h371e: o_data_a = 16'b1111110111101000;
            14'h371f: o_data_a = 16'b1110110010100000;
            14'h3720: o_data_a = 16'b1110001100001000;
            14'h3721: o_data_a = 16'b0000000000110011;
            14'h3722: o_data_a = 16'b1110110000010000;
            14'h3723: o_data_a = 16'b0000000000000000;
            14'h3724: o_data_a = 16'b1111110111101000;
            14'h3725: o_data_a = 16'b1110110010100000;
            14'h3726: o_data_a = 16'b1110001100001000;
            14'h3727: o_data_a = 16'b0000000000111111;
            14'h3728: o_data_a = 16'b1110110000010000;
            14'h3729: o_data_a = 16'b0000000000000000;
            14'h372a: o_data_a = 16'b1111110111101000;
            14'h372b: o_data_a = 16'b1110110010100000;
            14'h372c: o_data_a = 16'b1110001100001000;
            14'h372d: o_data_a = 16'b0000000000111011;
            14'h372e: o_data_a = 16'b1110110000010000;
            14'h372f: o_data_a = 16'b0000000000000000;
            14'h3730: o_data_a = 16'b1111110111101000;
            14'h3731: o_data_a = 16'b1110110010100000;
            14'h3732: o_data_a = 16'b1110001100001000;
            14'h3733: o_data_a = 16'b0000000000011110;
            14'h3734: o_data_a = 16'b1110110000010000;
            14'h3735: o_data_a = 16'b0000000000000000;
            14'h3736: o_data_a = 16'b1111110111101000;
            14'h3737: o_data_a = 16'b1110110010100000;
            14'h3738: o_data_a = 16'b1110001100001000;
            14'h3739: o_data_a = 16'b0000000000110000;
            14'h373a: o_data_a = 16'b1110110000010000;
            14'h373b: o_data_a = 16'b0000000000000000;
            14'h373c: o_data_a = 16'b1111110111101000;
            14'h373d: o_data_a = 16'b1110110010100000;
            14'h373e: o_data_a = 16'b1110001100001000;
            14'h373f: o_data_a = 16'b0000000000000000;
            14'h3740: o_data_a = 16'b1111110111001000;
            14'h3741: o_data_a = 16'b1111110010100000;
            14'h3742: o_data_a = 16'b1110101010001000;
            14'h3743: o_data_a = 16'b0000000000001100;
            14'h3744: o_data_a = 16'b1110110000010000;
            14'h3745: o_data_a = 16'b0000000000001101;
            14'h3746: o_data_a = 16'b1110001100001000;
            14'h3747: o_data_a = 16'b0100010110110011;
            14'h3748: o_data_a = 16'b1110110000010000;
            14'h3749: o_data_a = 16'b0000000000001110;
            14'h374a: o_data_a = 16'b1110001100001000;
            14'h374b: o_data_a = 16'b0011011101001111;
            14'h374c: o_data_a = 16'b1110110000010000;
            14'h374d: o_data_a = 16'b0000000001011111;
            14'h374e: o_data_a = 16'b1110101010000111;
            14'h374f: o_data_a = 16'b0000000000000000;
            14'h3750: o_data_a = 16'b1111110010101000;
            14'h3751: o_data_a = 16'b1111110000010000;
            14'h3752: o_data_a = 16'b0000000000000101;
            14'h3753: o_data_a = 16'b1110001100001000;
            14'h3754: o_data_a = 16'b0000000001010010;
            14'h3755: o_data_a = 16'b1110110000010000;
            14'h3756: o_data_a = 16'b0000000000000000;
            14'h3757: o_data_a = 16'b1111110111101000;
            14'h3758: o_data_a = 16'b1110110010100000;
            14'h3759: o_data_a = 16'b1110001100001000;
            14'h375a: o_data_a = 16'b0000000000011111;
            14'h375b: o_data_a = 16'b1110110000010000;
            14'h375c: o_data_a = 16'b0000000000000000;
            14'h375d: o_data_a = 16'b1111110111101000;
            14'h375e: o_data_a = 16'b1110110010100000;
            14'h375f: o_data_a = 16'b1110001100001000;
            14'h3760: o_data_a = 16'b0000000000110011;
            14'h3761: o_data_a = 16'b1110110000010000;
            14'h3762: o_data_a = 16'b0000000000000000;
            14'h3763: o_data_a = 16'b1111110111101000;
            14'h3764: o_data_a = 16'b1110110010100000;
            14'h3765: o_data_a = 16'b1110001100001000;
            14'h3766: o_data_a = 16'b0000000000110011;
            14'h3767: o_data_a = 16'b1110110000010000;
            14'h3768: o_data_a = 16'b0000000000000000;
            14'h3769: o_data_a = 16'b1111110111101000;
            14'h376a: o_data_a = 16'b1110110010100000;
            14'h376b: o_data_a = 16'b1110001100001000;
            14'h376c: o_data_a = 16'b0000000000110011;
            14'h376d: o_data_a = 16'b1110110000010000;
            14'h376e: o_data_a = 16'b0000000000000000;
            14'h376f: o_data_a = 16'b1111110111101000;
            14'h3770: o_data_a = 16'b1110110010100000;
            14'h3771: o_data_a = 16'b1110001100001000;
            14'h3772: o_data_a = 16'b0000000000011111;
            14'h3773: o_data_a = 16'b1110110000010000;
            14'h3774: o_data_a = 16'b0000000000000000;
            14'h3775: o_data_a = 16'b1111110111101000;
            14'h3776: o_data_a = 16'b1110110010100000;
            14'h3777: o_data_a = 16'b1110001100001000;
            14'h3778: o_data_a = 16'b0000000000011011;
            14'h3779: o_data_a = 16'b1110110000010000;
            14'h377a: o_data_a = 16'b0000000000000000;
            14'h377b: o_data_a = 16'b1111110111101000;
            14'h377c: o_data_a = 16'b1110110010100000;
            14'h377d: o_data_a = 16'b1110001100001000;
            14'h377e: o_data_a = 16'b0000000000110011;
            14'h377f: o_data_a = 16'b1110110000010000;
            14'h3780: o_data_a = 16'b0000000000000000;
            14'h3781: o_data_a = 16'b1111110111101000;
            14'h3782: o_data_a = 16'b1110110010100000;
            14'h3783: o_data_a = 16'b1110001100001000;
            14'h3784: o_data_a = 16'b0000000000110011;
            14'h3785: o_data_a = 16'b1110110000010000;
            14'h3786: o_data_a = 16'b0000000000000000;
            14'h3787: o_data_a = 16'b1111110111101000;
            14'h3788: o_data_a = 16'b1110110010100000;
            14'h3789: o_data_a = 16'b1110001100001000;
            14'h378a: o_data_a = 16'b0000000000110011;
            14'h378b: o_data_a = 16'b1110110000010000;
            14'h378c: o_data_a = 16'b0000000000000000;
            14'h378d: o_data_a = 16'b1111110111101000;
            14'h378e: o_data_a = 16'b1110110010100000;
            14'h378f: o_data_a = 16'b1110001100001000;
            14'h3790: o_data_a = 16'b0000000000000000;
            14'h3791: o_data_a = 16'b1111110111001000;
            14'h3792: o_data_a = 16'b1111110010100000;
            14'h3793: o_data_a = 16'b1110101010001000;
            14'h3794: o_data_a = 16'b0000000000000000;
            14'h3795: o_data_a = 16'b1111110111001000;
            14'h3796: o_data_a = 16'b1111110010100000;
            14'h3797: o_data_a = 16'b1110101010001000;
            14'h3798: o_data_a = 16'b0000000000001100;
            14'h3799: o_data_a = 16'b1110110000010000;
            14'h379a: o_data_a = 16'b0000000000001101;
            14'h379b: o_data_a = 16'b1110001100001000;
            14'h379c: o_data_a = 16'b0100010110110011;
            14'h379d: o_data_a = 16'b1110110000010000;
            14'h379e: o_data_a = 16'b0000000000001110;
            14'h379f: o_data_a = 16'b1110001100001000;
            14'h37a0: o_data_a = 16'b0011011110100100;
            14'h37a1: o_data_a = 16'b1110110000010000;
            14'h37a2: o_data_a = 16'b0000000001011111;
            14'h37a3: o_data_a = 16'b1110101010000111;
            14'h37a4: o_data_a = 16'b0000000000000000;
            14'h37a5: o_data_a = 16'b1111110010101000;
            14'h37a6: o_data_a = 16'b1111110000010000;
            14'h37a7: o_data_a = 16'b0000000000000101;
            14'h37a8: o_data_a = 16'b1110001100001000;
            14'h37a9: o_data_a = 16'b0000000001010011;
            14'h37aa: o_data_a = 16'b1110110000010000;
            14'h37ab: o_data_a = 16'b0000000000000000;
            14'h37ac: o_data_a = 16'b1111110111101000;
            14'h37ad: o_data_a = 16'b1110110010100000;
            14'h37ae: o_data_a = 16'b1110001100001000;
            14'h37af: o_data_a = 16'b0000000000011110;
            14'h37b0: o_data_a = 16'b1110110000010000;
            14'h37b1: o_data_a = 16'b0000000000000000;
            14'h37b2: o_data_a = 16'b1111110111101000;
            14'h37b3: o_data_a = 16'b1110110010100000;
            14'h37b4: o_data_a = 16'b1110001100001000;
            14'h37b5: o_data_a = 16'b0000000000110011;
            14'h37b6: o_data_a = 16'b1110110000010000;
            14'h37b7: o_data_a = 16'b0000000000000000;
            14'h37b8: o_data_a = 16'b1111110111101000;
            14'h37b9: o_data_a = 16'b1110110010100000;
            14'h37ba: o_data_a = 16'b1110001100001000;
            14'h37bb: o_data_a = 16'b0000000000110011;
            14'h37bc: o_data_a = 16'b1110110000010000;
            14'h37bd: o_data_a = 16'b0000000000000000;
            14'h37be: o_data_a = 16'b1111110111101000;
            14'h37bf: o_data_a = 16'b1110110010100000;
            14'h37c0: o_data_a = 16'b1110001100001000;
            14'h37c1: o_data_a = 16'b0000000000000110;
            14'h37c2: o_data_a = 16'b1110110000010000;
            14'h37c3: o_data_a = 16'b0000000000000000;
            14'h37c4: o_data_a = 16'b1111110111101000;
            14'h37c5: o_data_a = 16'b1110110010100000;
            14'h37c6: o_data_a = 16'b1110001100001000;
            14'h37c7: o_data_a = 16'b0000000000011100;
            14'h37c8: o_data_a = 16'b1110110000010000;
            14'h37c9: o_data_a = 16'b0000000000000000;
            14'h37ca: o_data_a = 16'b1111110111101000;
            14'h37cb: o_data_a = 16'b1110110010100000;
            14'h37cc: o_data_a = 16'b1110001100001000;
            14'h37cd: o_data_a = 16'b0000000000110000;
            14'h37ce: o_data_a = 16'b1110110000010000;
            14'h37cf: o_data_a = 16'b0000000000000000;
            14'h37d0: o_data_a = 16'b1111110111101000;
            14'h37d1: o_data_a = 16'b1110110010100000;
            14'h37d2: o_data_a = 16'b1110001100001000;
            14'h37d3: o_data_a = 16'b0000000000110011;
            14'h37d4: o_data_a = 16'b1110110000010000;
            14'h37d5: o_data_a = 16'b0000000000000000;
            14'h37d6: o_data_a = 16'b1111110111101000;
            14'h37d7: o_data_a = 16'b1110110010100000;
            14'h37d8: o_data_a = 16'b1110001100001000;
            14'h37d9: o_data_a = 16'b0000000000110011;
            14'h37da: o_data_a = 16'b1110110000010000;
            14'h37db: o_data_a = 16'b0000000000000000;
            14'h37dc: o_data_a = 16'b1111110111101000;
            14'h37dd: o_data_a = 16'b1110110010100000;
            14'h37de: o_data_a = 16'b1110001100001000;
            14'h37df: o_data_a = 16'b0000000000011110;
            14'h37e0: o_data_a = 16'b1110110000010000;
            14'h37e1: o_data_a = 16'b0000000000000000;
            14'h37e2: o_data_a = 16'b1111110111101000;
            14'h37e3: o_data_a = 16'b1110110010100000;
            14'h37e4: o_data_a = 16'b1110001100001000;
            14'h37e5: o_data_a = 16'b0000000000000000;
            14'h37e6: o_data_a = 16'b1111110111001000;
            14'h37e7: o_data_a = 16'b1111110010100000;
            14'h37e8: o_data_a = 16'b1110101010001000;
            14'h37e9: o_data_a = 16'b0000000000000000;
            14'h37ea: o_data_a = 16'b1111110111001000;
            14'h37eb: o_data_a = 16'b1111110010100000;
            14'h37ec: o_data_a = 16'b1110101010001000;
            14'h37ed: o_data_a = 16'b0000000000001100;
            14'h37ee: o_data_a = 16'b1110110000010000;
            14'h37ef: o_data_a = 16'b0000000000001101;
            14'h37f0: o_data_a = 16'b1110001100001000;
            14'h37f1: o_data_a = 16'b0100010110110011;
            14'h37f2: o_data_a = 16'b1110110000010000;
            14'h37f3: o_data_a = 16'b0000000000001110;
            14'h37f4: o_data_a = 16'b1110001100001000;
            14'h37f5: o_data_a = 16'b0011011111111001;
            14'h37f6: o_data_a = 16'b1110110000010000;
            14'h37f7: o_data_a = 16'b0000000001011111;
            14'h37f8: o_data_a = 16'b1110101010000111;
            14'h37f9: o_data_a = 16'b0000000000000000;
            14'h37fa: o_data_a = 16'b1111110010101000;
            14'h37fb: o_data_a = 16'b1111110000010000;
            14'h37fc: o_data_a = 16'b0000000000000101;
            14'h37fd: o_data_a = 16'b1110001100001000;
            14'h37fe: o_data_a = 16'b0000000001010100;
            14'h37ff: o_data_a = 16'b1110110000010000;
            14'h3800: o_data_a = 16'b0000000000000000;
            14'h3801: o_data_a = 16'b1111110111101000;
            14'h3802: o_data_a = 16'b1110110010100000;
            14'h3803: o_data_a = 16'b1110001100001000;
            14'h3804: o_data_a = 16'b0000000000111111;
            14'h3805: o_data_a = 16'b1110110000010000;
            14'h3806: o_data_a = 16'b0000000000000000;
            14'h3807: o_data_a = 16'b1111110111101000;
            14'h3808: o_data_a = 16'b1110110010100000;
            14'h3809: o_data_a = 16'b1110001100001000;
            14'h380a: o_data_a = 16'b0000000000111111;
            14'h380b: o_data_a = 16'b1110110000010000;
            14'h380c: o_data_a = 16'b0000000000000000;
            14'h380d: o_data_a = 16'b1111110111101000;
            14'h380e: o_data_a = 16'b1110110010100000;
            14'h380f: o_data_a = 16'b1110001100001000;
            14'h3810: o_data_a = 16'b0000000000101101;
            14'h3811: o_data_a = 16'b1110110000010000;
            14'h3812: o_data_a = 16'b0000000000000000;
            14'h3813: o_data_a = 16'b1111110111101000;
            14'h3814: o_data_a = 16'b1110110010100000;
            14'h3815: o_data_a = 16'b1110001100001000;
            14'h3816: o_data_a = 16'b0000000000001100;
            14'h3817: o_data_a = 16'b1110110000010000;
            14'h3818: o_data_a = 16'b0000000000000000;
            14'h3819: o_data_a = 16'b1111110111101000;
            14'h381a: o_data_a = 16'b1110110010100000;
            14'h381b: o_data_a = 16'b1110001100001000;
            14'h381c: o_data_a = 16'b0000000000001100;
            14'h381d: o_data_a = 16'b1110110000010000;
            14'h381e: o_data_a = 16'b0000000000000000;
            14'h381f: o_data_a = 16'b1111110111101000;
            14'h3820: o_data_a = 16'b1110110010100000;
            14'h3821: o_data_a = 16'b1110001100001000;
            14'h3822: o_data_a = 16'b0000000000001100;
            14'h3823: o_data_a = 16'b1110110000010000;
            14'h3824: o_data_a = 16'b0000000000000000;
            14'h3825: o_data_a = 16'b1111110111101000;
            14'h3826: o_data_a = 16'b1110110010100000;
            14'h3827: o_data_a = 16'b1110001100001000;
            14'h3828: o_data_a = 16'b0000000000001100;
            14'h3829: o_data_a = 16'b1110110000010000;
            14'h382a: o_data_a = 16'b0000000000000000;
            14'h382b: o_data_a = 16'b1111110111101000;
            14'h382c: o_data_a = 16'b1110110010100000;
            14'h382d: o_data_a = 16'b1110001100001000;
            14'h382e: o_data_a = 16'b0000000000001100;
            14'h382f: o_data_a = 16'b1110110000010000;
            14'h3830: o_data_a = 16'b0000000000000000;
            14'h3831: o_data_a = 16'b1111110111101000;
            14'h3832: o_data_a = 16'b1110110010100000;
            14'h3833: o_data_a = 16'b1110001100001000;
            14'h3834: o_data_a = 16'b0000000000011110;
            14'h3835: o_data_a = 16'b1110110000010000;
            14'h3836: o_data_a = 16'b0000000000000000;
            14'h3837: o_data_a = 16'b1111110111101000;
            14'h3838: o_data_a = 16'b1110110010100000;
            14'h3839: o_data_a = 16'b1110001100001000;
            14'h383a: o_data_a = 16'b0000000000000000;
            14'h383b: o_data_a = 16'b1111110111001000;
            14'h383c: o_data_a = 16'b1111110010100000;
            14'h383d: o_data_a = 16'b1110101010001000;
            14'h383e: o_data_a = 16'b0000000000000000;
            14'h383f: o_data_a = 16'b1111110111001000;
            14'h3840: o_data_a = 16'b1111110010100000;
            14'h3841: o_data_a = 16'b1110101010001000;
            14'h3842: o_data_a = 16'b0000000000001100;
            14'h3843: o_data_a = 16'b1110110000010000;
            14'h3844: o_data_a = 16'b0000000000001101;
            14'h3845: o_data_a = 16'b1110001100001000;
            14'h3846: o_data_a = 16'b0100010110110011;
            14'h3847: o_data_a = 16'b1110110000010000;
            14'h3848: o_data_a = 16'b0000000000001110;
            14'h3849: o_data_a = 16'b1110001100001000;
            14'h384a: o_data_a = 16'b0011100001001110;
            14'h384b: o_data_a = 16'b1110110000010000;
            14'h384c: o_data_a = 16'b0000000001011111;
            14'h384d: o_data_a = 16'b1110101010000111;
            14'h384e: o_data_a = 16'b0000000000000000;
            14'h384f: o_data_a = 16'b1111110010101000;
            14'h3850: o_data_a = 16'b1111110000010000;
            14'h3851: o_data_a = 16'b0000000000000101;
            14'h3852: o_data_a = 16'b1110001100001000;
            14'h3853: o_data_a = 16'b0000000001010101;
            14'h3854: o_data_a = 16'b1110110000010000;
            14'h3855: o_data_a = 16'b0000000000000000;
            14'h3856: o_data_a = 16'b1111110111101000;
            14'h3857: o_data_a = 16'b1110110010100000;
            14'h3858: o_data_a = 16'b1110001100001000;
            14'h3859: o_data_a = 16'b0000000000110011;
            14'h385a: o_data_a = 16'b1110110000010000;
            14'h385b: o_data_a = 16'b0000000000000000;
            14'h385c: o_data_a = 16'b1111110111101000;
            14'h385d: o_data_a = 16'b1110110010100000;
            14'h385e: o_data_a = 16'b1110001100001000;
            14'h385f: o_data_a = 16'b0000000000110011;
            14'h3860: o_data_a = 16'b1110110000010000;
            14'h3861: o_data_a = 16'b0000000000000000;
            14'h3862: o_data_a = 16'b1111110111101000;
            14'h3863: o_data_a = 16'b1110110010100000;
            14'h3864: o_data_a = 16'b1110001100001000;
            14'h3865: o_data_a = 16'b0000000000110011;
            14'h3866: o_data_a = 16'b1110110000010000;
            14'h3867: o_data_a = 16'b0000000000000000;
            14'h3868: o_data_a = 16'b1111110111101000;
            14'h3869: o_data_a = 16'b1110110010100000;
            14'h386a: o_data_a = 16'b1110001100001000;
            14'h386b: o_data_a = 16'b0000000000110011;
            14'h386c: o_data_a = 16'b1110110000010000;
            14'h386d: o_data_a = 16'b0000000000000000;
            14'h386e: o_data_a = 16'b1111110111101000;
            14'h386f: o_data_a = 16'b1110110010100000;
            14'h3870: o_data_a = 16'b1110001100001000;
            14'h3871: o_data_a = 16'b0000000000110011;
            14'h3872: o_data_a = 16'b1110110000010000;
            14'h3873: o_data_a = 16'b0000000000000000;
            14'h3874: o_data_a = 16'b1111110111101000;
            14'h3875: o_data_a = 16'b1110110010100000;
            14'h3876: o_data_a = 16'b1110001100001000;
            14'h3877: o_data_a = 16'b0000000000110011;
            14'h3878: o_data_a = 16'b1110110000010000;
            14'h3879: o_data_a = 16'b0000000000000000;
            14'h387a: o_data_a = 16'b1111110111101000;
            14'h387b: o_data_a = 16'b1110110010100000;
            14'h387c: o_data_a = 16'b1110001100001000;
            14'h387d: o_data_a = 16'b0000000000110011;
            14'h387e: o_data_a = 16'b1110110000010000;
            14'h387f: o_data_a = 16'b0000000000000000;
            14'h3880: o_data_a = 16'b1111110111101000;
            14'h3881: o_data_a = 16'b1110110010100000;
            14'h3882: o_data_a = 16'b1110001100001000;
            14'h3883: o_data_a = 16'b0000000000110011;
            14'h3884: o_data_a = 16'b1110110000010000;
            14'h3885: o_data_a = 16'b0000000000000000;
            14'h3886: o_data_a = 16'b1111110111101000;
            14'h3887: o_data_a = 16'b1110110010100000;
            14'h3888: o_data_a = 16'b1110001100001000;
            14'h3889: o_data_a = 16'b0000000000011110;
            14'h388a: o_data_a = 16'b1110110000010000;
            14'h388b: o_data_a = 16'b0000000000000000;
            14'h388c: o_data_a = 16'b1111110111101000;
            14'h388d: o_data_a = 16'b1110110010100000;
            14'h388e: o_data_a = 16'b1110001100001000;
            14'h388f: o_data_a = 16'b0000000000000000;
            14'h3890: o_data_a = 16'b1111110111001000;
            14'h3891: o_data_a = 16'b1111110010100000;
            14'h3892: o_data_a = 16'b1110101010001000;
            14'h3893: o_data_a = 16'b0000000000000000;
            14'h3894: o_data_a = 16'b1111110111001000;
            14'h3895: o_data_a = 16'b1111110010100000;
            14'h3896: o_data_a = 16'b1110101010001000;
            14'h3897: o_data_a = 16'b0000000000001100;
            14'h3898: o_data_a = 16'b1110110000010000;
            14'h3899: o_data_a = 16'b0000000000001101;
            14'h389a: o_data_a = 16'b1110001100001000;
            14'h389b: o_data_a = 16'b0100010110110011;
            14'h389c: o_data_a = 16'b1110110000010000;
            14'h389d: o_data_a = 16'b0000000000001110;
            14'h389e: o_data_a = 16'b1110001100001000;
            14'h389f: o_data_a = 16'b0011100010100011;
            14'h38a0: o_data_a = 16'b1110110000010000;
            14'h38a1: o_data_a = 16'b0000000001011111;
            14'h38a2: o_data_a = 16'b1110101010000111;
            14'h38a3: o_data_a = 16'b0000000000000000;
            14'h38a4: o_data_a = 16'b1111110010101000;
            14'h38a5: o_data_a = 16'b1111110000010000;
            14'h38a6: o_data_a = 16'b0000000000000101;
            14'h38a7: o_data_a = 16'b1110001100001000;
            14'h38a8: o_data_a = 16'b0000000001010110;
            14'h38a9: o_data_a = 16'b1110110000010000;
            14'h38aa: o_data_a = 16'b0000000000000000;
            14'h38ab: o_data_a = 16'b1111110111101000;
            14'h38ac: o_data_a = 16'b1110110010100000;
            14'h38ad: o_data_a = 16'b1110001100001000;
            14'h38ae: o_data_a = 16'b0000000000110011;
            14'h38af: o_data_a = 16'b1110110000010000;
            14'h38b0: o_data_a = 16'b0000000000000000;
            14'h38b1: o_data_a = 16'b1111110111101000;
            14'h38b2: o_data_a = 16'b1110110010100000;
            14'h38b3: o_data_a = 16'b1110001100001000;
            14'h38b4: o_data_a = 16'b0000000000110011;
            14'h38b5: o_data_a = 16'b1110110000010000;
            14'h38b6: o_data_a = 16'b0000000000000000;
            14'h38b7: o_data_a = 16'b1111110111101000;
            14'h38b8: o_data_a = 16'b1110110010100000;
            14'h38b9: o_data_a = 16'b1110001100001000;
            14'h38ba: o_data_a = 16'b0000000000110011;
            14'h38bb: o_data_a = 16'b1110110000010000;
            14'h38bc: o_data_a = 16'b0000000000000000;
            14'h38bd: o_data_a = 16'b1111110111101000;
            14'h38be: o_data_a = 16'b1110110010100000;
            14'h38bf: o_data_a = 16'b1110001100001000;
            14'h38c0: o_data_a = 16'b0000000000110011;
            14'h38c1: o_data_a = 16'b1110110000010000;
            14'h38c2: o_data_a = 16'b0000000000000000;
            14'h38c3: o_data_a = 16'b1111110111101000;
            14'h38c4: o_data_a = 16'b1110110010100000;
            14'h38c5: o_data_a = 16'b1110001100001000;
            14'h38c6: o_data_a = 16'b0000000000110011;
            14'h38c7: o_data_a = 16'b1110110000010000;
            14'h38c8: o_data_a = 16'b0000000000000000;
            14'h38c9: o_data_a = 16'b1111110111101000;
            14'h38ca: o_data_a = 16'b1110110010100000;
            14'h38cb: o_data_a = 16'b1110001100001000;
            14'h38cc: o_data_a = 16'b0000000000011110;
            14'h38cd: o_data_a = 16'b1110110000010000;
            14'h38ce: o_data_a = 16'b0000000000000000;
            14'h38cf: o_data_a = 16'b1111110111101000;
            14'h38d0: o_data_a = 16'b1110110010100000;
            14'h38d1: o_data_a = 16'b1110001100001000;
            14'h38d2: o_data_a = 16'b0000000000011110;
            14'h38d3: o_data_a = 16'b1110110000010000;
            14'h38d4: o_data_a = 16'b0000000000000000;
            14'h38d5: o_data_a = 16'b1111110111101000;
            14'h38d6: o_data_a = 16'b1110110010100000;
            14'h38d7: o_data_a = 16'b1110001100001000;
            14'h38d8: o_data_a = 16'b0000000000001100;
            14'h38d9: o_data_a = 16'b1110110000010000;
            14'h38da: o_data_a = 16'b0000000000000000;
            14'h38db: o_data_a = 16'b1111110111101000;
            14'h38dc: o_data_a = 16'b1110110010100000;
            14'h38dd: o_data_a = 16'b1110001100001000;
            14'h38de: o_data_a = 16'b0000000000001100;
            14'h38df: o_data_a = 16'b1110110000010000;
            14'h38e0: o_data_a = 16'b0000000000000000;
            14'h38e1: o_data_a = 16'b1111110111101000;
            14'h38e2: o_data_a = 16'b1110110010100000;
            14'h38e3: o_data_a = 16'b1110001100001000;
            14'h38e4: o_data_a = 16'b0000000000000000;
            14'h38e5: o_data_a = 16'b1111110111001000;
            14'h38e6: o_data_a = 16'b1111110010100000;
            14'h38e7: o_data_a = 16'b1110101010001000;
            14'h38e8: o_data_a = 16'b0000000000000000;
            14'h38e9: o_data_a = 16'b1111110111001000;
            14'h38ea: o_data_a = 16'b1111110010100000;
            14'h38eb: o_data_a = 16'b1110101010001000;
            14'h38ec: o_data_a = 16'b0000000000001100;
            14'h38ed: o_data_a = 16'b1110110000010000;
            14'h38ee: o_data_a = 16'b0000000000001101;
            14'h38ef: o_data_a = 16'b1110001100001000;
            14'h38f0: o_data_a = 16'b0100010110110011;
            14'h38f1: o_data_a = 16'b1110110000010000;
            14'h38f2: o_data_a = 16'b0000000000001110;
            14'h38f3: o_data_a = 16'b1110001100001000;
            14'h38f4: o_data_a = 16'b0011100011111000;
            14'h38f5: o_data_a = 16'b1110110000010000;
            14'h38f6: o_data_a = 16'b0000000001011111;
            14'h38f7: o_data_a = 16'b1110101010000111;
            14'h38f8: o_data_a = 16'b0000000000000000;
            14'h38f9: o_data_a = 16'b1111110010101000;
            14'h38fa: o_data_a = 16'b1111110000010000;
            14'h38fb: o_data_a = 16'b0000000000000101;
            14'h38fc: o_data_a = 16'b1110001100001000;
            14'h38fd: o_data_a = 16'b0000000001010111;
            14'h38fe: o_data_a = 16'b1110110000010000;
            14'h38ff: o_data_a = 16'b0000000000000000;
            14'h3900: o_data_a = 16'b1111110111101000;
            14'h3901: o_data_a = 16'b1110110010100000;
            14'h3902: o_data_a = 16'b1110001100001000;
            14'h3903: o_data_a = 16'b0000000000110011;
            14'h3904: o_data_a = 16'b1110110000010000;
            14'h3905: o_data_a = 16'b0000000000000000;
            14'h3906: o_data_a = 16'b1111110111101000;
            14'h3907: o_data_a = 16'b1110110010100000;
            14'h3908: o_data_a = 16'b1110001100001000;
            14'h3909: o_data_a = 16'b0000000000110011;
            14'h390a: o_data_a = 16'b1110110000010000;
            14'h390b: o_data_a = 16'b0000000000000000;
            14'h390c: o_data_a = 16'b1111110111101000;
            14'h390d: o_data_a = 16'b1110110010100000;
            14'h390e: o_data_a = 16'b1110001100001000;
            14'h390f: o_data_a = 16'b0000000000110011;
            14'h3910: o_data_a = 16'b1110110000010000;
            14'h3911: o_data_a = 16'b0000000000000000;
            14'h3912: o_data_a = 16'b1111110111101000;
            14'h3913: o_data_a = 16'b1110110010100000;
            14'h3914: o_data_a = 16'b1110001100001000;
            14'h3915: o_data_a = 16'b0000000000110011;
            14'h3916: o_data_a = 16'b1110110000010000;
            14'h3917: o_data_a = 16'b0000000000000000;
            14'h3918: o_data_a = 16'b1111110111101000;
            14'h3919: o_data_a = 16'b1110110010100000;
            14'h391a: o_data_a = 16'b1110001100001000;
            14'h391b: o_data_a = 16'b0000000000110011;
            14'h391c: o_data_a = 16'b1110110000010000;
            14'h391d: o_data_a = 16'b0000000000000000;
            14'h391e: o_data_a = 16'b1111110111101000;
            14'h391f: o_data_a = 16'b1110110010100000;
            14'h3920: o_data_a = 16'b1110001100001000;
            14'h3921: o_data_a = 16'b0000000000111111;
            14'h3922: o_data_a = 16'b1110110000010000;
            14'h3923: o_data_a = 16'b0000000000000000;
            14'h3924: o_data_a = 16'b1111110111101000;
            14'h3925: o_data_a = 16'b1110110010100000;
            14'h3926: o_data_a = 16'b1110001100001000;
            14'h3927: o_data_a = 16'b0000000000111111;
            14'h3928: o_data_a = 16'b1110110000010000;
            14'h3929: o_data_a = 16'b0000000000000000;
            14'h392a: o_data_a = 16'b1111110111101000;
            14'h392b: o_data_a = 16'b1110110010100000;
            14'h392c: o_data_a = 16'b1110001100001000;
            14'h392d: o_data_a = 16'b0000000000111111;
            14'h392e: o_data_a = 16'b1110110000010000;
            14'h392f: o_data_a = 16'b0000000000000000;
            14'h3930: o_data_a = 16'b1111110111101000;
            14'h3931: o_data_a = 16'b1110110010100000;
            14'h3932: o_data_a = 16'b1110001100001000;
            14'h3933: o_data_a = 16'b0000000000010010;
            14'h3934: o_data_a = 16'b1110110000010000;
            14'h3935: o_data_a = 16'b0000000000000000;
            14'h3936: o_data_a = 16'b1111110111101000;
            14'h3937: o_data_a = 16'b1110110010100000;
            14'h3938: o_data_a = 16'b1110001100001000;
            14'h3939: o_data_a = 16'b0000000000000000;
            14'h393a: o_data_a = 16'b1111110111001000;
            14'h393b: o_data_a = 16'b1111110010100000;
            14'h393c: o_data_a = 16'b1110101010001000;
            14'h393d: o_data_a = 16'b0000000000000000;
            14'h393e: o_data_a = 16'b1111110111001000;
            14'h393f: o_data_a = 16'b1111110010100000;
            14'h3940: o_data_a = 16'b1110101010001000;
            14'h3941: o_data_a = 16'b0000000000001100;
            14'h3942: o_data_a = 16'b1110110000010000;
            14'h3943: o_data_a = 16'b0000000000001101;
            14'h3944: o_data_a = 16'b1110001100001000;
            14'h3945: o_data_a = 16'b0100010110110011;
            14'h3946: o_data_a = 16'b1110110000010000;
            14'h3947: o_data_a = 16'b0000000000001110;
            14'h3948: o_data_a = 16'b1110001100001000;
            14'h3949: o_data_a = 16'b0011100101001101;
            14'h394a: o_data_a = 16'b1110110000010000;
            14'h394b: o_data_a = 16'b0000000001011111;
            14'h394c: o_data_a = 16'b1110101010000111;
            14'h394d: o_data_a = 16'b0000000000000000;
            14'h394e: o_data_a = 16'b1111110010101000;
            14'h394f: o_data_a = 16'b1111110000010000;
            14'h3950: o_data_a = 16'b0000000000000101;
            14'h3951: o_data_a = 16'b1110001100001000;
            14'h3952: o_data_a = 16'b0000000001011000;
            14'h3953: o_data_a = 16'b1110110000010000;
            14'h3954: o_data_a = 16'b0000000000000000;
            14'h3955: o_data_a = 16'b1111110111101000;
            14'h3956: o_data_a = 16'b1110110010100000;
            14'h3957: o_data_a = 16'b1110001100001000;
            14'h3958: o_data_a = 16'b0000000000110011;
            14'h3959: o_data_a = 16'b1110110000010000;
            14'h395a: o_data_a = 16'b0000000000000000;
            14'h395b: o_data_a = 16'b1111110111101000;
            14'h395c: o_data_a = 16'b1110110010100000;
            14'h395d: o_data_a = 16'b1110001100001000;
            14'h395e: o_data_a = 16'b0000000000110011;
            14'h395f: o_data_a = 16'b1110110000010000;
            14'h3960: o_data_a = 16'b0000000000000000;
            14'h3961: o_data_a = 16'b1111110111101000;
            14'h3962: o_data_a = 16'b1110110010100000;
            14'h3963: o_data_a = 16'b1110001100001000;
            14'h3964: o_data_a = 16'b0000000000011110;
            14'h3965: o_data_a = 16'b1110110000010000;
            14'h3966: o_data_a = 16'b0000000000000000;
            14'h3967: o_data_a = 16'b1111110111101000;
            14'h3968: o_data_a = 16'b1110110010100000;
            14'h3969: o_data_a = 16'b1110001100001000;
            14'h396a: o_data_a = 16'b0000000000011110;
            14'h396b: o_data_a = 16'b1110110000010000;
            14'h396c: o_data_a = 16'b0000000000000000;
            14'h396d: o_data_a = 16'b1111110111101000;
            14'h396e: o_data_a = 16'b1110110010100000;
            14'h396f: o_data_a = 16'b1110001100001000;
            14'h3970: o_data_a = 16'b0000000000001100;
            14'h3971: o_data_a = 16'b1110110000010000;
            14'h3972: o_data_a = 16'b0000000000000000;
            14'h3973: o_data_a = 16'b1111110111101000;
            14'h3974: o_data_a = 16'b1110110010100000;
            14'h3975: o_data_a = 16'b1110001100001000;
            14'h3976: o_data_a = 16'b0000000000011110;
            14'h3977: o_data_a = 16'b1110110000010000;
            14'h3978: o_data_a = 16'b0000000000000000;
            14'h3979: o_data_a = 16'b1111110111101000;
            14'h397a: o_data_a = 16'b1110110010100000;
            14'h397b: o_data_a = 16'b1110001100001000;
            14'h397c: o_data_a = 16'b0000000000011110;
            14'h397d: o_data_a = 16'b1110110000010000;
            14'h397e: o_data_a = 16'b0000000000000000;
            14'h397f: o_data_a = 16'b1111110111101000;
            14'h3980: o_data_a = 16'b1110110010100000;
            14'h3981: o_data_a = 16'b1110001100001000;
            14'h3982: o_data_a = 16'b0000000000110011;
            14'h3983: o_data_a = 16'b1110110000010000;
            14'h3984: o_data_a = 16'b0000000000000000;
            14'h3985: o_data_a = 16'b1111110111101000;
            14'h3986: o_data_a = 16'b1110110010100000;
            14'h3987: o_data_a = 16'b1110001100001000;
            14'h3988: o_data_a = 16'b0000000000110011;
            14'h3989: o_data_a = 16'b1110110000010000;
            14'h398a: o_data_a = 16'b0000000000000000;
            14'h398b: o_data_a = 16'b1111110111101000;
            14'h398c: o_data_a = 16'b1110110010100000;
            14'h398d: o_data_a = 16'b1110001100001000;
            14'h398e: o_data_a = 16'b0000000000000000;
            14'h398f: o_data_a = 16'b1111110111001000;
            14'h3990: o_data_a = 16'b1111110010100000;
            14'h3991: o_data_a = 16'b1110101010001000;
            14'h3992: o_data_a = 16'b0000000000000000;
            14'h3993: o_data_a = 16'b1111110111001000;
            14'h3994: o_data_a = 16'b1111110010100000;
            14'h3995: o_data_a = 16'b1110101010001000;
            14'h3996: o_data_a = 16'b0000000000001100;
            14'h3997: o_data_a = 16'b1110110000010000;
            14'h3998: o_data_a = 16'b0000000000001101;
            14'h3999: o_data_a = 16'b1110001100001000;
            14'h399a: o_data_a = 16'b0100010110110011;
            14'h399b: o_data_a = 16'b1110110000010000;
            14'h399c: o_data_a = 16'b0000000000001110;
            14'h399d: o_data_a = 16'b1110001100001000;
            14'h399e: o_data_a = 16'b0011100110100010;
            14'h399f: o_data_a = 16'b1110110000010000;
            14'h39a0: o_data_a = 16'b0000000001011111;
            14'h39a1: o_data_a = 16'b1110101010000111;
            14'h39a2: o_data_a = 16'b0000000000000000;
            14'h39a3: o_data_a = 16'b1111110010101000;
            14'h39a4: o_data_a = 16'b1111110000010000;
            14'h39a5: o_data_a = 16'b0000000000000101;
            14'h39a6: o_data_a = 16'b1110001100001000;
            14'h39a7: o_data_a = 16'b0000000001011001;
            14'h39a8: o_data_a = 16'b1110110000010000;
            14'h39a9: o_data_a = 16'b0000000000000000;
            14'h39aa: o_data_a = 16'b1111110111101000;
            14'h39ab: o_data_a = 16'b1110110010100000;
            14'h39ac: o_data_a = 16'b1110001100001000;
            14'h39ad: o_data_a = 16'b0000000000110011;
            14'h39ae: o_data_a = 16'b1110110000010000;
            14'h39af: o_data_a = 16'b0000000000000000;
            14'h39b0: o_data_a = 16'b1111110111101000;
            14'h39b1: o_data_a = 16'b1110110010100000;
            14'h39b2: o_data_a = 16'b1110001100001000;
            14'h39b3: o_data_a = 16'b0000000000110011;
            14'h39b4: o_data_a = 16'b1110110000010000;
            14'h39b5: o_data_a = 16'b0000000000000000;
            14'h39b6: o_data_a = 16'b1111110111101000;
            14'h39b7: o_data_a = 16'b1110110010100000;
            14'h39b8: o_data_a = 16'b1110001100001000;
            14'h39b9: o_data_a = 16'b0000000000110011;
            14'h39ba: o_data_a = 16'b1110110000010000;
            14'h39bb: o_data_a = 16'b0000000000000000;
            14'h39bc: o_data_a = 16'b1111110111101000;
            14'h39bd: o_data_a = 16'b1110110010100000;
            14'h39be: o_data_a = 16'b1110001100001000;
            14'h39bf: o_data_a = 16'b0000000000110011;
            14'h39c0: o_data_a = 16'b1110110000010000;
            14'h39c1: o_data_a = 16'b0000000000000000;
            14'h39c2: o_data_a = 16'b1111110111101000;
            14'h39c3: o_data_a = 16'b1110110010100000;
            14'h39c4: o_data_a = 16'b1110001100001000;
            14'h39c5: o_data_a = 16'b0000000000011110;
            14'h39c6: o_data_a = 16'b1110110000010000;
            14'h39c7: o_data_a = 16'b0000000000000000;
            14'h39c8: o_data_a = 16'b1111110111101000;
            14'h39c9: o_data_a = 16'b1110110010100000;
            14'h39ca: o_data_a = 16'b1110001100001000;
            14'h39cb: o_data_a = 16'b0000000000001100;
            14'h39cc: o_data_a = 16'b1110110000010000;
            14'h39cd: o_data_a = 16'b0000000000000000;
            14'h39ce: o_data_a = 16'b1111110111101000;
            14'h39cf: o_data_a = 16'b1110110010100000;
            14'h39d0: o_data_a = 16'b1110001100001000;
            14'h39d1: o_data_a = 16'b0000000000001100;
            14'h39d2: o_data_a = 16'b1110110000010000;
            14'h39d3: o_data_a = 16'b0000000000000000;
            14'h39d4: o_data_a = 16'b1111110111101000;
            14'h39d5: o_data_a = 16'b1110110010100000;
            14'h39d6: o_data_a = 16'b1110001100001000;
            14'h39d7: o_data_a = 16'b0000000000001100;
            14'h39d8: o_data_a = 16'b1110110000010000;
            14'h39d9: o_data_a = 16'b0000000000000000;
            14'h39da: o_data_a = 16'b1111110111101000;
            14'h39db: o_data_a = 16'b1110110010100000;
            14'h39dc: o_data_a = 16'b1110001100001000;
            14'h39dd: o_data_a = 16'b0000000000011110;
            14'h39de: o_data_a = 16'b1110110000010000;
            14'h39df: o_data_a = 16'b0000000000000000;
            14'h39e0: o_data_a = 16'b1111110111101000;
            14'h39e1: o_data_a = 16'b1110110010100000;
            14'h39e2: o_data_a = 16'b1110001100001000;
            14'h39e3: o_data_a = 16'b0000000000000000;
            14'h39e4: o_data_a = 16'b1111110111001000;
            14'h39e5: o_data_a = 16'b1111110010100000;
            14'h39e6: o_data_a = 16'b1110101010001000;
            14'h39e7: o_data_a = 16'b0000000000000000;
            14'h39e8: o_data_a = 16'b1111110111001000;
            14'h39e9: o_data_a = 16'b1111110010100000;
            14'h39ea: o_data_a = 16'b1110101010001000;
            14'h39eb: o_data_a = 16'b0000000000001100;
            14'h39ec: o_data_a = 16'b1110110000010000;
            14'h39ed: o_data_a = 16'b0000000000001101;
            14'h39ee: o_data_a = 16'b1110001100001000;
            14'h39ef: o_data_a = 16'b0100010110110011;
            14'h39f0: o_data_a = 16'b1110110000010000;
            14'h39f1: o_data_a = 16'b0000000000001110;
            14'h39f2: o_data_a = 16'b1110001100001000;
            14'h39f3: o_data_a = 16'b0011100111110111;
            14'h39f4: o_data_a = 16'b1110110000010000;
            14'h39f5: o_data_a = 16'b0000000001011111;
            14'h39f6: o_data_a = 16'b1110101010000111;
            14'h39f7: o_data_a = 16'b0000000000000000;
            14'h39f8: o_data_a = 16'b1111110010101000;
            14'h39f9: o_data_a = 16'b1111110000010000;
            14'h39fa: o_data_a = 16'b0000000000000101;
            14'h39fb: o_data_a = 16'b1110001100001000;
            14'h39fc: o_data_a = 16'b0000000001011010;
            14'h39fd: o_data_a = 16'b1110110000010000;
            14'h39fe: o_data_a = 16'b0000000000000000;
            14'h39ff: o_data_a = 16'b1111110111101000;
            14'h3a00: o_data_a = 16'b1110110010100000;
            14'h3a01: o_data_a = 16'b1110001100001000;
            14'h3a02: o_data_a = 16'b0000000000111111;
            14'h3a03: o_data_a = 16'b1110110000010000;
            14'h3a04: o_data_a = 16'b0000000000000000;
            14'h3a05: o_data_a = 16'b1111110111101000;
            14'h3a06: o_data_a = 16'b1110110010100000;
            14'h3a07: o_data_a = 16'b1110001100001000;
            14'h3a08: o_data_a = 16'b0000000000110011;
            14'h3a09: o_data_a = 16'b1110110000010000;
            14'h3a0a: o_data_a = 16'b0000000000000000;
            14'h3a0b: o_data_a = 16'b1111110111101000;
            14'h3a0c: o_data_a = 16'b1110110010100000;
            14'h3a0d: o_data_a = 16'b1110001100001000;
            14'h3a0e: o_data_a = 16'b0000000000110001;
            14'h3a0f: o_data_a = 16'b1110110000010000;
            14'h3a10: o_data_a = 16'b0000000000000000;
            14'h3a11: o_data_a = 16'b1111110111101000;
            14'h3a12: o_data_a = 16'b1110110010100000;
            14'h3a13: o_data_a = 16'b1110001100001000;
            14'h3a14: o_data_a = 16'b0000000000011000;
            14'h3a15: o_data_a = 16'b1110110000010000;
            14'h3a16: o_data_a = 16'b0000000000000000;
            14'h3a17: o_data_a = 16'b1111110111101000;
            14'h3a18: o_data_a = 16'b1110110010100000;
            14'h3a19: o_data_a = 16'b1110001100001000;
            14'h3a1a: o_data_a = 16'b0000000000001100;
            14'h3a1b: o_data_a = 16'b1110110000010000;
            14'h3a1c: o_data_a = 16'b0000000000000000;
            14'h3a1d: o_data_a = 16'b1111110111101000;
            14'h3a1e: o_data_a = 16'b1110110010100000;
            14'h3a1f: o_data_a = 16'b1110001100001000;
            14'h3a20: o_data_a = 16'b0000000000000110;
            14'h3a21: o_data_a = 16'b1110110000010000;
            14'h3a22: o_data_a = 16'b0000000000000000;
            14'h3a23: o_data_a = 16'b1111110111101000;
            14'h3a24: o_data_a = 16'b1110110010100000;
            14'h3a25: o_data_a = 16'b1110001100001000;
            14'h3a26: o_data_a = 16'b0000000000100011;
            14'h3a27: o_data_a = 16'b1110110000010000;
            14'h3a28: o_data_a = 16'b0000000000000000;
            14'h3a29: o_data_a = 16'b1111110111101000;
            14'h3a2a: o_data_a = 16'b1110110010100000;
            14'h3a2b: o_data_a = 16'b1110001100001000;
            14'h3a2c: o_data_a = 16'b0000000000110011;
            14'h3a2d: o_data_a = 16'b1110110000010000;
            14'h3a2e: o_data_a = 16'b0000000000000000;
            14'h3a2f: o_data_a = 16'b1111110111101000;
            14'h3a30: o_data_a = 16'b1110110010100000;
            14'h3a31: o_data_a = 16'b1110001100001000;
            14'h3a32: o_data_a = 16'b0000000000111111;
            14'h3a33: o_data_a = 16'b1110110000010000;
            14'h3a34: o_data_a = 16'b0000000000000000;
            14'h3a35: o_data_a = 16'b1111110111101000;
            14'h3a36: o_data_a = 16'b1110110010100000;
            14'h3a37: o_data_a = 16'b1110001100001000;
            14'h3a38: o_data_a = 16'b0000000000000000;
            14'h3a39: o_data_a = 16'b1111110111001000;
            14'h3a3a: o_data_a = 16'b1111110010100000;
            14'h3a3b: o_data_a = 16'b1110101010001000;
            14'h3a3c: o_data_a = 16'b0000000000000000;
            14'h3a3d: o_data_a = 16'b1111110111001000;
            14'h3a3e: o_data_a = 16'b1111110010100000;
            14'h3a3f: o_data_a = 16'b1110101010001000;
            14'h3a40: o_data_a = 16'b0000000000001100;
            14'h3a41: o_data_a = 16'b1110110000010000;
            14'h3a42: o_data_a = 16'b0000000000001101;
            14'h3a43: o_data_a = 16'b1110001100001000;
            14'h3a44: o_data_a = 16'b0100010110110011;
            14'h3a45: o_data_a = 16'b1110110000010000;
            14'h3a46: o_data_a = 16'b0000000000001110;
            14'h3a47: o_data_a = 16'b1110001100001000;
            14'h3a48: o_data_a = 16'b0011101001001100;
            14'h3a49: o_data_a = 16'b1110110000010000;
            14'h3a4a: o_data_a = 16'b0000000001011111;
            14'h3a4b: o_data_a = 16'b1110101010000111;
            14'h3a4c: o_data_a = 16'b0000000000000000;
            14'h3a4d: o_data_a = 16'b1111110010101000;
            14'h3a4e: o_data_a = 16'b1111110000010000;
            14'h3a4f: o_data_a = 16'b0000000000000101;
            14'h3a50: o_data_a = 16'b1110001100001000;
            14'h3a51: o_data_a = 16'b0000000001011011;
            14'h3a52: o_data_a = 16'b1110110000010000;
            14'h3a53: o_data_a = 16'b0000000000000000;
            14'h3a54: o_data_a = 16'b1111110111101000;
            14'h3a55: o_data_a = 16'b1110110010100000;
            14'h3a56: o_data_a = 16'b1110001100001000;
            14'h3a57: o_data_a = 16'b0000000000011110;
            14'h3a58: o_data_a = 16'b1110110000010000;
            14'h3a59: o_data_a = 16'b0000000000000000;
            14'h3a5a: o_data_a = 16'b1111110111101000;
            14'h3a5b: o_data_a = 16'b1110110010100000;
            14'h3a5c: o_data_a = 16'b1110001100001000;
            14'h3a5d: o_data_a = 16'b0000000000000110;
            14'h3a5e: o_data_a = 16'b1110110000010000;
            14'h3a5f: o_data_a = 16'b0000000000000000;
            14'h3a60: o_data_a = 16'b1111110111101000;
            14'h3a61: o_data_a = 16'b1110110010100000;
            14'h3a62: o_data_a = 16'b1110001100001000;
            14'h3a63: o_data_a = 16'b0000000000000110;
            14'h3a64: o_data_a = 16'b1110110000010000;
            14'h3a65: o_data_a = 16'b0000000000000000;
            14'h3a66: o_data_a = 16'b1111110111101000;
            14'h3a67: o_data_a = 16'b1110110010100000;
            14'h3a68: o_data_a = 16'b1110001100001000;
            14'h3a69: o_data_a = 16'b0000000000000110;
            14'h3a6a: o_data_a = 16'b1110110000010000;
            14'h3a6b: o_data_a = 16'b0000000000000000;
            14'h3a6c: o_data_a = 16'b1111110111101000;
            14'h3a6d: o_data_a = 16'b1110110010100000;
            14'h3a6e: o_data_a = 16'b1110001100001000;
            14'h3a6f: o_data_a = 16'b0000000000000110;
            14'h3a70: o_data_a = 16'b1110110000010000;
            14'h3a71: o_data_a = 16'b0000000000000000;
            14'h3a72: o_data_a = 16'b1111110111101000;
            14'h3a73: o_data_a = 16'b1110110010100000;
            14'h3a74: o_data_a = 16'b1110001100001000;
            14'h3a75: o_data_a = 16'b0000000000000110;
            14'h3a76: o_data_a = 16'b1110110000010000;
            14'h3a77: o_data_a = 16'b0000000000000000;
            14'h3a78: o_data_a = 16'b1111110111101000;
            14'h3a79: o_data_a = 16'b1110110010100000;
            14'h3a7a: o_data_a = 16'b1110001100001000;
            14'h3a7b: o_data_a = 16'b0000000000000110;
            14'h3a7c: o_data_a = 16'b1110110000010000;
            14'h3a7d: o_data_a = 16'b0000000000000000;
            14'h3a7e: o_data_a = 16'b1111110111101000;
            14'h3a7f: o_data_a = 16'b1110110010100000;
            14'h3a80: o_data_a = 16'b1110001100001000;
            14'h3a81: o_data_a = 16'b0000000000000110;
            14'h3a82: o_data_a = 16'b1110110000010000;
            14'h3a83: o_data_a = 16'b0000000000000000;
            14'h3a84: o_data_a = 16'b1111110111101000;
            14'h3a85: o_data_a = 16'b1110110010100000;
            14'h3a86: o_data_a = 16'b1110001100001000;
            14'h3a87: o_data_a = 16'b0000000000011110;
            14'h3a88: o_data_a = 16'b1110110000010000;
            14'h3a89: o_data_a = 16'b0000000000000000;
            14'h3a8a: o_data_a = 16'b1111110111101000;
            14'h3a8b: o_data_a = 16'b1110110010100000;
            14'h3a8c: o_data_a = 16'b1110001100001000;
            14'h3a8d: o_data_a = 16'b0000000000000000;
            14'h3a8e: o_data_a = 16'b1111110111001000;
            14'h3a8f: o_data_a = 16'b1111110010100000;
            14'h3a90: o_data_a = 16'b1110101010001000;
            14'h3a91: o_data_a = 16'b0000000000000000;
            14'h3a92: o_data_a = 16'b1111110111001000;
            14'h3a93: o_data_a = 16'b1111110010100000;
            14'h3a94: o_data_a = 16'b1110101010001000;
            14'h3a95: o_data_a = 16'b0000000000001100;
            14'h3a96: o_data_a = 16'b1110110000010000;
            14'h3a97: o_data_a = 16'b0000000000001101;
            14'h3a98: o_data_a = 16'b1110001100001000;
            14'h3a99: o_data_a = 16'b0100010110110011;
            14'h3a9a: o_data_a = 16'b1110110000010000;
            14'h3a9b: o_data_a = 16'b0000000000001110;
            14'h3a9c: o_data_a = 16'b1110001100001000;
            14'h3a9d: o_data_a = 16'b0011101010100001;
            14'h3a9e: o_data_a = 16'b1110110000010000;
            14'h3a9f: o_data_a = 16'b0000000001011111;
            14'h3aa0: o_data_a = 16'b1110101010000111;
            14'h3aa1: o_data_a = 16'b0000000000000000;
            14'h3aa2: o_data_a = 16'b1111110010101000;
            14'h3aa3: o_data_a = 16'b1111110000010000;
            14'h3aa4: o_data_a = 16'b0000000000000101;
            14'h3aa5: o_data_a = 16'b1110001100001000;
            14'h3aa6: o_data_a = 16'b0000000001011100;
            14'h3aa7: o_data_a = 16'b1110110000010000;
            14'h3aa8: o_data_a = 16'b0000000000000000;
            14'h3aa9: o_data_a = 16'b1111110111101000;
            14'h3aaa: o_data_a = 16'b1110110010100000;
            14'h3aab: o_data_a = 16'b1110001100001000;
            14'h3aac: o_data_a = 16'b0000000000000000;
            14'h3aad: o_data_a = 16'b1111110111001000;
            14'h3aae: o_data_a = 16'b1111110010100000;
            14'h3aaf: o_data_a = 16'b1110101010001000;
            14'h3ab0: o_data_a = 16'b0000000000000000;
            14'h3ab1: o_data_a = 16'b1111110111001000;
            14'h3ab2: o_data_a = 16'b1111110010100000;
            14'h3ab3: o_data_a = 16'b1110101010001000;
            14'h3ab4: o_data_a = 16'b0000000000000000;
            14'h3ab5: o_data_a = 16'b1111110111001000;
            14'h3ab6: o_data_a = 16'b1111110010100000;
            14'h3ab7: o_data_a = 16'b1110111111001000;
            14'h3ab8: o_data_a = 16'b0000000000000011;
            14'h3ab9: o_data_a = 16'b1110110000010000;
            14'h3aba: o_data_a = 16'b0000000000000000;
            14'h3abb: o_data_a = 16'b1111110111101000;
            14'h3abc: o_data_a = 16'b1110110010100000;
            14'h3abd: o_data_a = 16'b1110001100001000;
            14'h3abe: o_data_a = 16'b0000000000000110;
            14'h3abf: o_data_a = 16'b1110110000010000;
            14'h3ac0: o_data_a = 16'b0000000000000000;
            14'h3ac1: o_data_a = 16'b1111110111101000;
            14'h3ac2: o_data_a = 16'b1110110010100000;
            14'h3ac3: o_data_a = 16'b1110001100001000;
            14'h3ac4: o_data_a = 16'b0000000000001100;
            14'h3ac5: o_data_a = 16'b1110110000010000;
            14'h3ac6: o_data_a = 16'b0000000000000000;
            14'h3ac7: o_data_a = 16'b1111110111101000;
            14'h3ac8: o_data_a = 16'b1110110010100000;
            14'h3ac9: o_data_a = 16'b1110001100001000;
            14'h3aca: o_data_a = 16'b0000000000011000;
            14'h3acb: o_data_a = 16'b1110110000010000;
            14'h3acc: o_data_a = 16'b0000000000000000;
            14'h3acd: o_data_a = 16'b1111110111101000;
            14'h3ace: o_data_a = 16'b1110110010100000;
            14'h3acf: o_data_a = 16'b1110001100001000;
            14'h3ad0: o_data_a = 16'b0000000000110000;
            14'h3ad1: o_data_a = 16'b1110110000010000;
            14'h3ad2: o_data_a = 16'b0000000000000000;
            14'h3ad3: o_data_a = 16'b1111110111101000;
            14'h3ad4: o_data_a = 16'b1110110010100000;
            14'h3ad5: o_data_a = 16'b1110001100001000;
            14'h3ad6: o_data_a = 16'b0000000000100000;
            14'h3ad7: o_data_a = 16'b1110110000010000;
            14'h3ad8: o_data_a = 16'b0000000000000000;
            14'h3ad9: o_data_a = 16'b1111110111101000;
            14'h3ada: o_data_a = 16'b1110110010100000;
            14'h3adb: o_data_a = 16'b1110001100001000;
            14'h3adc: o_data_a = 16'b0000000000000000;
            14'h3add: o_data_a = 16'b1111110111001000;
            14'h3ade: o_data_a = 16'b1111110010100000;
            14'h3adf: o_data_a = 16'b1110101010001000;
            14'h3ae0: o_data_a = 16'b0000000000000000;
            14'h3ae1: o_data_a = 16'b1111110111001000;
            14'h3ae2: o_data_a = 16'b1111110010100000;
            14'h3ae3: o_data_a = 16'b1110101010001000;
            14'h3ae4: o_data_a = 16'b0000000000001100;
            14'h3ae5: o_data_a = 16'b1110110000010000;
            14'h3ae6: o_data_a = 16'b0000000000001101;
            14'h3ae7: o_data_a = 16'b1110001100001000;
            14'h3ae8: o_data_a = 16'b0100010110110011;
            14'h3ae9: o_data_a = 16'b1110110000010000;
            14'h3aea: o_data_a = 16'b0000000000001110;
            14'h3aeb: o_data_a = 16'b1110001100001000;
            14'h3aec: o_data_a = 16'b0011101011110000;
            14'h3aed: o_data_a = 16'b1110110000010000;
            14'h3aee: o_data_a = 16'b0000000001011111;
            14'h3aef: o_data_a = 16'b1110101010000111;
            14'h3af0: o_data_a = 16'b0000000000000000;
            14'h3af1: o_data_a = 16'b1111110010101000;
            14'h3af2: o_data_a = 16'b1111110000010000;
            14'h3af3: o_data_a = 16'b0000000000000101;
            14'h3af4: o_data_a = 16'b1110001100001000;
            14'h3af5: o_data_a = 16'b0000000001011101;
            14'h3af6: o_data_a = 16'b1110110000010000;
            14'h3af7: o_data_a = 16'b0000000000000000;
            14'h3af8: o_data_a = 16'b1111110111101000;
            14'h3af9: o_data_a = 16'b1110110010100000;
            14'h3afa: o_data_a = 16'b1110001100001000;
            14'h3afb: o_data_a = 16'b0000000000011110;
            14'h3afc: o_data_a = 16'b1110110000010000;
            14'h3afd: o_data_a = 16'b0000000000000000;
            14'h3afe: o_data_a = 16'b1111110111101000;
            14'h3aff: o_data_a = 16'b1110110010100000;
            14'h3b00: o_data_a = 16'b1110001100001000;
            14'h3b01: o_data_a = 16'b0000000000011000;
            14'h3b02: o_data_a = 16'b1110110000010000;
            14'h3b03: o_data_a = 16'b0000000000000000;
            14'h3b04: o_data_a = 16'b1111110111101000;
            14'h3b05: o_data_a = 16'b1110110010100000;
            14'h3b06: o_data_a = 16'b1110001100001000;
            14'h3b07: o_data_a = 16'b0000000000011000;
            14'h3b08: o_data_a = 16'b1110110000010000;
            14'h3b09: o_data_a = 16'b0000000000000000;
            14'h3b0a: o_data_a = 16'b1111110111101000;
            14'h3b0b: o_data_a = 16'b1110110010100000;
            14'h3b0c: o_data_a = 16'b1110001100001000;
            14'h3b0d: o_data_a = 16'b0000000000011000;
            14'h3b0e: o_data_a = 16'b1110110000010000;
            14'h3b0f: o_data_a = 16'b0000000000000000;
            14'h3b10: o_data_a = 16'b1111110111101000;
            14'h3b11: o_data_a = 16'b1110110010100000;
            14'h3b12: o_data_a = 16'b1110001100001000;
            14'h3b13: o_data_a = 16'b0000000000011000;
            14'h3b14: o_data_a = 16'b1110110000010000;
            14'h3b15: o_data_a = 16'b0000000000000000;
            14'h3b16: o_data_a = 16'b1111110111101000;
            14'h3b17: o_data_a = 16'b1110110010100000;
            14'h3b18: o_data_a = 16'b1110001100001000;
            14'h3b19: o_data_a = 16'b0000000000011000;
            14'h3b1a: o_data_a = 16'b1110110000010000;
            14'h3b1b: o_data_a = 16'b0000000000000000;
            14'h3b1c: o_data_a = 16'b1111110111101000;
            14'h3b1d: o_data_a = 16'b1110110010100000;
            14'h3b1e: o_data_a = 16'b1110001100001000;
            14'h3b1f: o_data_a = 16'b0000000000011000;
            14'h3b20: o_data_a = 16'b1110110000010000;
            14'h3b21: o_data_a = 16'b0000000000000000;
            14'h3b22: o_data_a = 16'b1111110111101000;
            14'h3b23: o_data_a = 16'b1110110010100000;
            14'h3b24: o_data_a = 16'b1110001100001000;
            14'h3b25: o_data_a = 16'b0000000000011000;
            14'h3b26: o_data_a = 16'b1110110000010000;
            14'h3b27: o_data_a = 16'b0000000000000000;
            14'h3b28: o_data_a = 16'b1111110111101000;
            14'h3b29: o_data_a = 16'b1110110010100000;
            14'h3b2a: o_data_a = 16'b1110001100001000;
            14'h3b2b: o_data_a = 16'b0000000000011110;
            14'h3b2c: o_data_a = 16'b1110110000010000;
            14'h3b2d: o_data_a = 16'b0000000000000000;
            14'h3b2e: o_data_a = 16'b1111110111101000;
            14'h3b2f: o_data_a = 16'b1110110010100000;
            14'h3b30: o_data_a = 16'b1110001100001000;
            14'h3b31: o_data_a = 16'b0000000000000000;
            14'h3b32: o_data_a = 16'b1111110111001000;
            14'h3b33: o_data_a = 16'b1111110010100000;
            14'h3b34: o_data_a = 16'b1110101010001000;
            14'h3b35: o_data_a = 16'b0000000000000000;
            14'h3b36: o_data_a = 16'b1111110111001000;
            14'h3b37: o_data_a = 16'b1111110010100000;
            14'h3b38: o_data_a = 16'b1110101010001000;
            14'h3b39: o_data_a = 16'b0000000000001100;
            14'h3b3a: o_data_a = 16'b1110110000010000;
            14'h3b3b: o_data_a = 16'b0000000000001101;
            14'h3b3c: o_data_a = 16'b1110001100001000;
            14'h3b3d: o_data_a = 16'b0100010110110011;
            14'h3b3e: o_data_a = 16'b1110110000010000;
            14'h3b3f: o_data_a = 16'b0000000000001110;
            14'h3b40: o_data_a = 16'b1110001100001000;
            14'h3b41: o_data_a = 16'b0011101101000101;
            14'h3b42: o_data_a = 16'b1110110000010000;
            14'h3b43: o_data_a = 16'b0000000001011111;
            14'h3b44: o_data_a = 16'b1110101010000111;
            14'h3b45: o_data_a = 16'b0000000000000000;
            14'h3b46: o_data_a = 16'b1111110010101000;
            14'h3b47: o_data_a = 16'b1111110000010000;
            14'h3b48: o_data_a = 16'b0000000000000101;
            14'h3b49: o_data_a = 16'b1110001100001000;
            14'h3b4a: o_data_a = 16'b0000000001011110;
            14'h3b4b: o_data_a = 16'b1110110000010000;
            14'h3b4c: o_data_a = 16'b0000000000000000;
            14'h3b4d: o_data_a = 16'b1111110111101000;
            14'h3b4e: o_data_a = 16'b1110110010100000;
            14'h3b4f: o_data_a = 16'b1110001100001000;
            14'h3b50: o_data_a = 16'b0000000000001000;
            14'h3b51: o_data_a = 16'b1110110000010000;
            14'h3b52: o_data_a = 16'b0000000000000000;
            14'h3b53: o_data_a = 16'b1111110111101000;
            14'h3b54: o_data_a = 16'b1110110010100000;
            14'h3b55: o_data_a = 16'b1110001100001000;
            14'h3b56: o_data_a = 16'b0000000000011100;
            14'h3b57: o_data_a = 16'b1110110000010000;
            14'h3b58: o_data_a = 16'b0000000000000000;
            14'h3b59: o_data_a = 16'b1111110111101000;
            14'h3b5a: o_data_a = 16'b1110110010100000;
            14'h3b5b: o_data_a = 16'b1110001100001000;
            14'h3b5c: o_data_a = 16'b0000000000110110;
            14'h3b5d: o_data_a = 16'b1110110000010000;
            14'h3b5e: o_data_a = 16'b0000000000000000;
            14'h3b5f: o_data_a = 16'b1111110111101000;
            14'h3b60: o_data_a = 16'b1110110010100000;
            14'h3b61: o_data_a = 16'b1110001100001000;
            14'h3b62: o_data_a = 16'b0000000000000000;
            14'h3b63: o_data_a = 16'b1111110111001000;
            14'h3b64: o_data_a = 16'b1111110010100000;
            14'h3b65: o_data_a = 16'b1110101010001000;
            14'h3b66: o_data_a = 16'b0000000000000000;
            14'h3b67: o_data_a = 16'b1111110111001000;
            14'h3b68: o_data_a = 16'b1111110010100000;
            14'h3b69: o_data_a = 16'b1110101010001000;
            14'h3b6a: o_data_a = 16'b0000000000000000;
            14'h3b6b: o_data_a = 16'b1111110111001000;
            14'h3b6c: o_data_a = 16'b1111110010100000;
            14'h3b6d: o_data_a = 16'b1110101010001000;
            14'h3b6e: o_data_a = 16'b0000000000000000;
            14'h3b6f: o_data_a = 16'b1111110111001000;
            14'h3b70: o_data_a = 16'b1111110010100000;
            14'h3b71: o_data_a = 16'b1110101010001000;
            14'h3b72: o_data_a = 16'b0000000000000000;
            14'h3b73: o_data_a = 16'b1111110111001000;
            14'h3b74: o_data_a = 16'b1111110010100000;
            14'h3b75: o_data_a = 16'b1110101010001000;
            14'h3b76: o_data_a = 16'b0000000000000000;
            14'h3b77: o_data_a = 16'b1111110111001000;
            14'h3b78: o_data_a = 16'b1111110010100000;
            14'h3b79: o_data_a = 16'b1110101010001000;
            14'h3b7a: o_data_a = 16'b0000000000000000;
            14'h3b7b: o_data_a = 16'b1111110111001000;
            14'h3b7c: o_data_a = 16'b1111110010100000;
            14'h3b7d: o_data_a = 16'b1110101010001000;
            14'h3b7e: o_data_a = 16'b0000000000000000;
            14'h3b7f: o_data_a = 16'b1111110111001000;
            14'h3b80: o_data_a = 16'b1111110010100000;
            14'h3b81: o_data_a = 16'b1110101010001000;
            14'h3b82: o_data_a = 16'b0000000000001100;
            14'h3b83: o_data_a = 16'b1110110000010000;
            14'h3b84: o_data_a = 16'b0000000000001101;
            14'h3b85: o_data_a = 16'b1110001100001000;
            14'h3b86: o_data_a = 16'b0100010110110011;
            14'h3b87: o_data_a = 16'b1110110000010000;
            14'h3b88: o_data_a = 16'b0000000000001110;
            14'h3b89: o_data_a = 16'b1110001100001000;
            14'h3b8a: o_data_a = 16'b0011101110001110;
            14'h3b8b: o_data_a = 16'b1110110000010000;
            14'h3b8c: o_data_a = 16'b0000000001011111;
            14'h3b8d: o_data_a = 16'b1110101010000111;
            14'h3b8e: o_data_a = 16'b0000000000000000;
            14'h3b8f: o_data_a = 16'b1111110010101000;
            14'h3b90: o_data_a = 16'b1111110000010000;
            14'h3b91: o_data_a = 16'b0000000000000101;
            14'h3b92: o_data_a = 16'b1110001100001000;
            14'h3b93: o_data_a = 16'b0000000001011111;
            14'h3b94: o_data_a = 16'b1110110000010000;
            14'h3b95: o_data_a = 16'b0000000000000000;
            14'h3b96: o_data_a = 16'b1111110111101000;
            14'h3b97: o_data_a = 16'b1110110010100000;
            14'h3b98: o_data_a = 16'b1110001100001000;
            14'h3b99: o_data_a = 16'b0000000000000000;
            14'h3b9a: o_data_a = 16'b1111110111001000;
            14'h3b9b: o_data_a = 16'b1111110010100000;
            14'h3b9c: o_data_a = 16'b1110101010001000;
            14'h3b9d: o_data_a = 16'b0000000000000000;
            14'h3b9e: o_data_a = 16'b1111110111001000;
            14'h3b9f: o_data_a = 16'b1111110010100000;
            14'h3ba0: o_data_a = 16'b1110101010001000;
            14'h3ba1: o_data_a = 16'b0000000000000000;
            14'h3ba2: o_data_a = 16'b1111110111001000;
            14'h3ba3: o_data_a = 16'b1111110010100000;
            14'h3ba4: o_data_a = 16'b1110101010001000;
            14'h3ba5: o_data_a = 16'b0000000000000000;
            14'h3ba6: o_data_a = 16'b1111110111001000;
            14'h3ba7: o_data_a = 16'b1111110010100000;
            14'h3ba8: o_data_a = 16'b1110101010001000;
            14'h3ba9: o_data_a = 16'b0000000000000000;
            14'h3baa: o_data_a = 16'b1111110111001000;
            14'h3bab: o_data_a = 16'b1111110010100000;
            14'h3bac: o_data_a = 16'b1110101010001000;
            14'h3bad: o_data_a = 16'b0000000000000000;
            14'h3bae: o_data_a = 16'b1111110111001000;
            14'h3baf: o_data_a = 16'b1111110010100000;
            14'h3bb0: o_data_a = 16'b1110101010001000;
            14'h3bb1: o_data_a = 16'b0000000000000000;
            14'h3bb2: o_data_a = 16'b1111110111001000;
            14'h3bb3: o_data_a = 16'b1111110010100000;
            14'h3bb4: o_data_a = 16'b1110101010001000;
            14'h3bb5: o_data_a = 16'b0000000000000000;
            14'h3bb6: o_data_a = 16'b1111110111001000;
            14'h3bb7: o_data_a = 16'b1111110010100000;
            14'h3bb8: o_data_a = 16'b1110101010001000;
            14'h3bb9: o_data_a = 16'b0000000000000000;
            14'h3bba: o_data_a = 16'b1111110111001000;
            14'h3bbb: o_data_a = 16'b1111110010100000;
            14'h3bbc: o_data_a = 16'b1110101010001000;
            14'h3bbd: o_data_a = 16'b0000000000111111;
            14'h3bbe: o_data_a = 16'b1110110000010000;
            14'h3bbf: o_data_a = 16'b0000000000000000;
            14'h3bc0: o_data_a = 16'b1111110111101000;
            14'h3bc1: o_data_a = 16'b1110110010100000;
            14'h3bc2: o_data_a = 16'b1110001100001000;
            14'h3bc3: o_data_a = 16'b0000000000000000;
            14'h3bc4: o_data_a = 16'b1111110111001000;
            14'h3bc5: o_data_a = 16'b1111110010100000;
            14'h3bc6: o_data_a = 16'b1110101010001000;
            14'h3bc7: o_data_a = 16'b0000000000001100;
            14'h3bc8: o_data_a = 16'b1110110000010000;
            14'h3bc9: o_data_a = 16'b0000000000001101;
            14'h3bca: o_data_a = 16'b1110001100001000;
            14'h3bcb: o_data_a = 16'b0100010110110011;
            14'h3bcc: o_data_a = 16'b1110110000010000;
            14'h3bcd: o_data_a = 16'b0000000000001110;
            14'h3bce: o_data_a = 16'b1110001100001000;
            14'h3bcf: o_data_a = 16'b0011101111010011;
            14'h3bd0: o_data_a = 16'b1110110000010000;
            14'h3bd1: o_data_a = 16'b0000000001011111;
            14'h3bd2: o_data_a = 16'b1110101010000111;
            14'h3bd3: o_data_a = 16'b0000000000000000;
            14'h3bd4: o_data_a = 16'b1111110010101000;
            14'h3bd5: o_data_a = 16'b1111110000010000;
            14'h3bd6: o_data_a = 16'b0000000000000101;
            14'h3bd7: o_data_a = 16'b1110001100001000;
            14'h3bd8: o_data_a = 16'b0000000001100000;
            14'h3bd9: o_data_a = 16'b1110110000010000;
            14'h3bda: o_data_a = 16'b0000000000000000;
            14'h3bdb: o_data_a = 16'b1111110111101000;
            14'h3bdc: o_data_a = 16'b1110110010100000;
            14'h3bdd: o_data_a = 16'b1110001100001000;
            14'h3bde: o_data_a = 16'b0000000000000110;
            14'h3bdf: o_data_a = 16'b1110110000010000;
            14'h3be0: o_data_a = 16'b0000000000000000;
            14'h3be1: o_data_a = 16'b1111110111101000;
            14'h3be2: o_data_a = 16'b1110110010100000;
            14'h3be3: o_data_a = 16'b1110001100001000;
            14'h3be4: o_data_a = 16'b0000000000001100;
            14'h3be5: o_data_a = 16'b1110110000010000;
            14'h3be6: o_data_a = 16'b0000000000000000;
            14'h3be7: o_data_a = 16'b1111110111101000;
            14'h3be8: o_data_a = 16'b1110110010100000;
            14'h3be9: o_data_a = 16'b1110001100001000;
            14'h3bea: o_data_a = 16'b0000000000011000;
            14'h3beb: o_data_a = 16'b1110110000010000;
            14'h3bec: o_data_a = 16'b0000000000000000;
            14'h3bed: o_data_a = 16'b1111110111101000;
            14'h3bee: o_data_a = 16'b1110110010100000;
            14'h3bef: o_data_a = 16'b1110001100001000;
            14'h3bf0: o_data_a = 16'b0000000000000000;
            14'h3bf1: o_data_a = 16'b1111110111001000;
            14'h3bf2: o_data_a = 16'b1111110010100000;
            14'h3bf3: o_data_a = 16'b1110101010001000;
            14'h3bf4: o_data_a = 16'b0000000000000000;
            14'h3bf5: o_data_a = 16'b1111110111001000;
            14'h3bf6: o_data_a = 16'b1111110010100000;
            14'h3bf7: o_data_a = 16'b1110101010001000;
            14'h3bf8: o_data_a = 16'b0000000000000000;
            14'h3bf9: o_data_a = 16'b1111110111001000;
            14'h3bfa: o_data_a = 16'b1111110010100000;
            14'h3bfb: o_data_a = 16'b1110101010001000;
            14'h3bfc: o_data_a = 16'b0000000000000000;
            14'h3bfd: o_data_a = 16'b1111110111001000;
            14'h3bfe: o_data_a = 16'b1111110010100000;
            14'h3bff: o_data_a = 16'b1110101010001000;
            14'h3c00: o_data_a = 16'b0000000000000000;
            14'h3c01: o_data_a = 16'b1111110111001000;
            14'h3c02: o_data_a = 16'b1111110010100000;
            14'h3c03: o_data_a = 16'b1110101010001000;
            14'h3c04: o_data_a = 16'b0000000000000000;
            14'h3c05: o_data_a = 16'b1111110111001000;
            14'h3c06: o_data_a = 16'b1111110010100000;
            14'h3c07: o_data_a = 16'b1110101010001000;
            14'h3c08: o_data_a = 16'b0000000000000000;
            14'h3c09: o_data_a = 16'b1111110111001000;
            14'h3c0a: o_data_a = 16'b1111110010100000;
            14'h3c0b: o_data_a = 16'b1110101010001000;
            14'h3c0c: o_data_a = 16'b0000000000000000;
            14'h3c0d: o_data_a = 16'b1111110111001000;
            14'h3c0e: o_data_a = 16'b1111110010100000;
            14'h3c0f: o_data_a = 16'b1110101010001000;
            14'h3c10: o_data_a = 16'b0000000000001100;
            14'h3c11: o_data_a = 16'b1110110000010000;
            14'h3c12: o_data_a = 16'b0000000000001101;
            14'h3c13: o_data_a = 16'b1110001100001000;
            14'h3c14: o_data_a = 16'b0100010110110011;
            14'h3c15: o_data_a = 16'b1110110000010000;
            14'h3c16: o_data_a = 16'b0000000000001110;
            14'h3c17: o_data_a = 16'b1110001100001000;
            14'h3c18: o_data_a = 16'b0011110000011100;
            14'h3c19: o_data_a = 16'b1110110000010000;
            14'h3c1a: o_data_a = 16'b0000000001011111;
            14'h3c1b: o_data_a = 16'b1110101010000111;
            14'h3c1c: o_data_a = 16'b0000000000000000;
            14'h3c1d: o_data_a = 16'b1111110010101000;
            14'h3c1e: o_data_a = 16'b1111110000010000;
            14'h3c1f: o_data_a = 16'b0000000000000101;
            14'h3c20: o_data_a = 16'b1110001100001000;
            14'h3c21: o_data_a = 16'b0000000001100001;
            14'h3c22: o_data_a = 16'b1110110000010000;
            14'h3c23: o_data_a = 16'b0000000000000000;
            14'h3c24: o_data_a = 16'b1111110111101000;
            14'h3c25: o_data_a = 16'b1110110010100000;
            14'h3c26: o_data_a = 16'b1110001100001000;
            14'h3c27: o_data_a = 16'b0000000000000000;
            14'h3c28: o_data_a = 16'b1111110111001000;
            14'h3c29: o_data_a = 16'b1111110010100000;
            14'h3c2a: o_data_a = 16'b1110101010001000;
            14'h3c2b: o_data_a = 16'b0000000000000000;
            14'h3c2c: o_data_a = 16'b1111110111001000;
            14'h3c2d: o_data_a = 16'b1111110010100000;
            14'h3c2e: o_data_a = 16'b1110101010001000;
            14'h3c2f: o_data_a = 16'b0000000000000000;
            14'h3c30: o_data_a = 16'b1111110111001000;
            14'h3c31: o_data_a = 16'b1111110010100000;
            14'h3c32: o_data_a = 16'b1110101010001000;
            14'h3c33: o_data_a = 16'b0000000000001110;
            14'h3c34: o_data_a = 16'b1110110000010000;
            14'h3c35: o_data_a = 16'b0000000000000000;
            14'h3c36: o_data_a = 16'b1111110111101000;
            14'h3c37: o_data_a = 16'b1110110010100000;
            14'h3c38: o_data_a = 16'b1110001100001000;
            14'h3c39: o_data_a = 16'b0000000000011000;
            14'h3c3a: o_data_a = 16'b1110110000010000;
            14'h3c3b: o_data_a = 16'b0000000000000000;
            14'h3c3c: o_data_a = 16'b1111110111101000;
            14'h3c3d: o_data_a = 16'b1110110010100000;
            14'h3c3e: o_data_a = 16'b1110001100001000;
            14'h3c3f: o_data_a = 16'b0000000000011110;
            14'h3c40: o_data_a = 16'b1110110000010000;
            14'h3c41: o_data_a = 16'b0000000000000000;
            14'h3c42: o_data_a = 16'b1111110111101000;
            14'h3c43: o_data_a = 16'b1110110010100000;
            14'h3c44: o_data_a = 16'b1110001100001000;
            14'h3c45: o_data_a = 16'b0000000000011011;
            14'h3c46: o_data_a = 16'b1110110000010000;
            14'h3c47: o_data_a = 16'b0000000000000000;
            14'h3c48: o_data_a = 16'b1111110111101000;
            14'h3c49: o_data_a = 16'b1110110010100000;
            14'h3c4a: o_data_a = 16'b1110001100001000;
            14'h3c4b: o_data_a = 16'b0000000000011011;
            14'h3c4c: o_data_a = 16'b1110110000010000;
            14'h3c4d: o_data_a = 16'b0000000000000000;
            14'h3c4e: o_data_a = 16'b1111110111101000;
            14'h3c4f: o_data_a = 16'b1110110010100000;
            14'h3c50: o_data_a = 16'b1110001100001000;
            14'h3c51: o_data_a = 16'b0000000000110110;
            14'h3c52: o_data_a = 16'b1110110000010000;
            14'h3c53: o_data_a = 16'b0000000000000000;
            14'h3c54: o_data_a = 16'b1111110111101000;
            14'h3c55: o_data_a = 16'b1110110010100000;
            14'h3c56: o_data_a = 16'b1110001100001000;
            14'h3c57: o_data_a = 16'b0000000000000000;
            14'h3c58: o_data_a = 16'b1111110111001000;
            14'h3c59: o_data_a = 16'b1111110010100000;
            14'h3c5a: o_data_a = 16'b1110101010001000;
            14'h3c5b: o_data_a = 16'b0000000000000000;
            14'h3c5c: o_data_a = 16'b1111110111001000;
            14'h3c5d: o_data_a = 16'b1111110010100000;
            14'h3c5e: o_data_a = 16'b1110101010001000;
            14'h3c5f: o_data_a = 16'b0000000000001100;
            14'h3c60: o_data_a = 16'b1110110000010000;
            14'h3c61: o_data_a = 16'b0000000000001101;
            14'h3c62: o_data_a = 16'b1110001100001000;
            14'h3c63: o_data_a = 16'b0100010110110011;
            14'h3c64: o_data_a = 16'b1110110000010000;
            14'h3c65: o_data_a = 16'b0000000000001110;
            14'h3c66: o_data_a = 16'b1110001100001000;
            14'h3c67: o_data_a = 16'b0011110001101011;
            14'h3c68: o_data_a = 16'b1110110000010000;
            14'h3c69: o_data_a = 16'b0000000001011111;
            14'h3c6a: o_data_a = 16'b1110101010000111;
            14'h3c6b: o_data_a = 16'b0000000000000000;
            14'h3c6c: o_data_a = 16'b1111110010101000;
            14'h3c6d: o_data_a = 16'b1111110000010000;
            14'h3c6e: o_data_a = 16'b0000000000000101;
            14'h3c6f: o_data_a = 16'b1110001100001000;
            14'h3c70: o_data_a = 16'b0000000001100010;
            14'h3c71: o_data_a = 16'b1110110000010000;
            14'h3c72: o_data_a = 16'b0000000000000000;
            14'h3c73: o_data_a = 16'b1111110111101000;
            14'h3c74: o_data_a = 16'b1110110010100000;
            14'h3c75: o_data_a = 16'b1110001100001000;
            14'h3c76: o_data_a = 16'b0000000000000011;
            14'h3c77: o_data_a = 16'b1110110000010000;
            14'h3c78: o_data_a = 16'b0000000000000000;
            14'h3c79: o_data_a = 16'b1111110111101000;
            14'h3c7a: o_data_a = 16'b1110110010100000;
            14'h3c7b: o_data_a = 16'b1110001100001000;
            14'h3c7c: o_data_a = 16'b0000000000000011;
            14'h3c7d: o_data_a = 16'b1110110000010000;
            14'h3c7e: o_data_a = 16'b0000000000000000;
            14'h3c7f: o_data_a = 16'b1111110111101000;
            14'h3c80: o_data_a = 16'b1110110010100000;
            14'h3c81: o_data_a = 16'b1110001100001000;
            14'h3c82: o_data_a = 16'b0000000000000011;
            14'h3c83: o_data_a = 16'b1110110000010000;
            14'h3c84: o_data_a = 16'b0000000000000000;
            14'h3c85: o_data_a = 16'b1111110111101000;
            14'h3c86: o_data_a = 16'b1110110010100000;
            14'h3c87: o_data_a = 16'b1110001100001000;
            14'h3c88: o_data_a = 16'b0000000000001111;
            14'h3c89: o_data_a = 16'b1110110000010000;
            14'h3c8a: o_data_a = 16'b0000000000000000;
            14'h3c8b: o_data_a = 16'b1111110111101000;
            14'h3c8c: o_data_a = 16'b1110110010100000;
            14'h3c8d: o_data_a = 16'b1110001100001000;
            14'h3c8e: o_data_a = 16'b0000000000011011;
            14'h3c8f: o_data_a = 16'b1110110000010000;
            14'h3c90: o_data_a = 16'b0000000000000000;
            14'h3c91: o_data_a = 16'b1111110111101000;
            14'h3c92: o_data_a = 16'b1110110010100000;
            14'h3c93: o_data_a = 16'b1110001100001000;
            14'h3c94: o_data_a = 16'b0000000000110011;
            14'h3c95: o_data_a = 16'b1110110000010000;
            14'h3c96: o_data_a = 16'b0000000000000000;
            14'h3c97: o_data_a = 16'b1111110111101000;
            14'h3c98: o_data_a = 16'b1110110010100000;
            14'h3c99: o_data_a = 16'b1110001100001000;
            14'h3c9a: o_data_a = 16'b0000000000110011;
            14'h3c9b: o_data_a = 16'b1110110000010000;
            14'h3c9c: o_data_a = 16'b0000000000000000;
            14'h3c9d: o_data_a = 16'b1111110111101000;
            14'h3c9e: o_data_a = 16'b1110110010100000;
            14'h3c9f: o_data_a = 16'b1110001100001000;
            14'h3ca0: o_data_a = 16'b0000000000110011;
            14'h3ca1: o_data_a = 16'b1110110000010000;
            14'h3ca2: o_data_a = 16'b0000000000000000;
            14'h3ca3: o_data_a = 16'b1111110111101000;
            14'h3ca4: o_data_a = 16'b1110110010100000;
            14'h3ca5: o_data_a = 16'b1110001100001000;
            14'h3ca6: o_data_a = 16'b0000000000011110;
            14'h3ca7: o_data_a = 16'b1110110000010000;
            14'h3ca8: o_data_a = 16'b0000000000000000;
            14'h3ca9: o_data_a = 16'b1111110111101000;
            14'h3caa: o_data_a = 16'b1110110010100000;
            14'h3cab: o_data_a = 16'b1110001100001000;
            14'h3cac: o_data_a = 16'b0000000000000000;
            14'h3cad: o_data_a = 16'b1111110111001000;
            14'h3cae: o_data_a = 16'b1111110010100000;
            14'h3caf: o_data_a = 16'b1110101010001000;
            14'h3cb0: o_data_a = 16'b0000000000000000;
            14'h3cb1: o_data_a = 16'b1111110111001000;
            14'h3cb2: o_data_a = 16'b1111110010100000;
            14'h3cb3: o_data_a = 16'b1110101010001000;
            14'h3cb4: o_data_a = 16'b0000000000001100;
            14'h3cb5: o_data_a = 16'b1110110000010000;
            14'h3cb6: o_data_a = 16'b0000000000001101;
            14'h3cb7: o_data_a = 16'b1110001100001000;
            14'h3cb8: o_data_a = 16'b0100010110110011;
            14'h3cb9: o_data_a = 16'b1110110000010000;
            14'h3cba: o_data_a = 16'b0000000000001110;
            14'h3cbb: o_data_a = 16'b1110001100001000;
            14'h3cbc: o_data_a = 16'b0011110011000000;
            14'h3cbd: o_data_a = 16'b1110110000010000;
            14'h3cbe: o_data_a = 16'b0000000001011111;
            14'h3cbf: o_data_a = 16'b1110101010000111;
            14'h3cc0: o_data_a = 16'b0000000000000000;
            14'h3cc1: o_data_a = 16'b1111110010101000;
            14'h3cc2: o_data_a = 16'b1111110000010000;
            14'h3cc3: o_data_a = 16'b0000000000000101;
            14'h3cc4: o_data_a = 16'b1110001100001000;
            14'h3cc5: o_data_a = 16'b0000000001100011;
            14'h3cc6: o_data_a = 16'b1110110000010000;
            14'h3cc7: o_data_a = 16'b0000000000000000;
            14'h3cc8: o_data_a = 16'b1111110111101000;
            14'h3cc9: o_data_a = 16'b1110110010100000;
            14'h3cca: o_data_a = 16'b1110001100001000;
            14'h3ccb: o_data_a = 16'b0000000000000000;
            14'h3ccc: o_data_a = 16'b1111110111001000;
            14'h3ccd: o_data_a = 16'b1111110010100000;
            14'h3cce: o_data_a = 16'b1110101010001000;
            14'h3ccf: o_data_a = 16'b0000000000000000;
            14'h3cd0: o_data_a = 16'b1111110111001000;
            14'h3cd1: o_data_a = 16'b1111110010100000;
            14'h3cd2: o_data_a = 16'b1110101010001000;
            14'h3cd3: o_data_a = 16'b0000000000000000;
            14'h3cd4: o_data_a = 16'b1111110111001000;
            14'h3cd5: o_data_a = 16'b1111110010100000;
            14'h3cd6: o_data_a = 16'b1110101010001000;
            14'h3cd7: o_data_a = 16'b0000000000011110;
            14'h3cd8: o_data_a = 16'b1110110000010000;
            14'h3cd9: o_data_a = 16'b0000000000000000;
            14'h3cda: o_data_a = 16'b1111110111101000;
            14'h3cdb: o_data_a = 16'b1110110010100000;
            14'h3cdc: o_data_a = 16'b1110001100001000;
            14'h3cdd: o_data_a = 16'b0000000000110011;
            14'h3cde: o_data_a = 16'b1110110000010000;
            14'h3cdf: o_data_a = 16'b0000000000000000;
            14'h3ce0: o_data_a = 16'b1111110111101000;
            14'h3ce1: o_data_a = 16'b1110110010100000;
            14'h3ce2: o_data_a = 16'b1110001100001000;
            14'h3ce3: o_data_a = 16'b0000000000000011;
            14'h3ce4: o_data_a = 16'b1110110000010000;
            14'h3ce5: o_data_a = 16'b0000000000000000;
            14'h3ce6: o_data_a = 16'b1111110111101000;
            14'h3ce7: o_data_a = 16'b1110110010100000;
            14'h3ce8: o_data_a = 16'b1110001100001000;
            14'h3ce9: o_data_a = 16'b0000000000000011;
            14'h3cea: o_data_a = 16'b1110110000010000;
            14'h3ceb: o_data_a = 16'b0000000000000000;
            14'h3cec: o_data_a = 16'b1111110111101000;
            14'h3ced: o_data_a = 16'b1110110010100000;
            14'h3cee: o_data_a = 16'b1110001100001000;
            14'h3cef: o_data_a = 16'b0000000000110011;
            14'h3cf0: o_data_a = 16'b1110110000010000;
            14'h3cf1: o_data_a = 16'b0000000000000000;
            14'h3cf2: o_data_a = 16'b1111110111101000;
            14'h3cf3: o_data_a = 16'b1110110010100000;
            14'h3cf4: o_data_a = 16'b1110001100001000;
            14'h3cf5: o_data_a = 16'b0000000000011110;
            14'h3cf6: o_data_a = 16'b1110110000010000;
            14'h3cf7: o_data_a = 16'b0000000000000000;
            14'h3cf8: o_data_a = 16'b1111110111101000;
            14'h3cf9: o_data_a = 16'b1110110010100000;
            14'h3cfa: o_data_a = 16'b1110001100001000;
            14'h3cfb: o_data_a = 16'b0000000000000000;
            14'h3cfc: o_data_a = 16'b1111110111001000;
            14'h3cfd: o_data_a = 16'b1111110010100000;
            14'h3cfe: o_data_a = 16'b1110101010001000;
            14'h3cff: o_data_a = 16'b0000000000000000;
            14'h3d00: o_data_a = 16'b1111110111001000;
            14'h3d01: o_data_a = 16'b1111110010100000;
            14'h3d02: o_data_a = 16'b1110101010001000;
            14'h3d03: o_data_a = 16'b0000000000001100;
            14'h3d04: o_data_a = 16'b1110110000010000;
            14'h3d05: o_data_a = 16'b0000000000001101;
            14'h3d06: o_data_a = 16'b1110001100001000;
            14'h3d07: o_data_a = 16'b0100010110110011;
            14'h3d08: o_data_a = 16'b1110110000010000;
            14'h3d09: o_data_a = 16'b0000000000001110;
            14'h3d0a: o_data_a = 16'b1110001100001000;
            14'h3d0b: o_data_a = 16'b0011110100001111;
            14'h3d0c: o_data_a = 16'b1110110000010000;
            14'h3d0d: o_data_a = 16'b0000000001011111;
            14'h3d0e: o_data_a = 16'b1110101010000111;
            14'h3d0f: o_data_a = 16'b0000000000000000;
            14'h3d10: o_data_a = 16'b1111110010101000;
            14'h3d11: o_data_a = 16'b1111110000010000;
            14'h3d12: o_data_a = 16'b0000000000000101;
            14'h3d13: o_data_a = 16'b1110001100001000;
            14'h3d14: o_data_a = 16'b0000000001100100;
            14'h3d15: o_data_a = 16'b1110110000010000;
            14'h3d16: o_data_a = 16'b0000000000000000;
            14'h3d17: o_data_a = 16'b1111110111101000;
            14'h3d18: o_data_a = 16'b1110110010100000;
            14'h3d19: o_data_a = 16'b1110001100001000;
            14'h3d1a: o_data_a = 16'b0000000000110000;
            14'h3d1b: o_data_a = 16'b1110110000010000;
            14'h3d1c: o_data_a = 16'b0000000000000000;
            14'h3d1d: o_data_a = 16'b1111110111101000;
            14'h3d1e: o_data_a = 16'b1110110010100000;
            14'h3d1f: o_data_a = 16'b1110001100001000;
            14'h3d20: o_data_a = 16'b0000000000110000;
            14'h3d21: o_data_a = 16'b1110110000010000;
            14'h3d22: o_data_a = 16'b0000000000000000;
            14'h3d23: o_data_a = 16'b1111110111101000;
            14'h3d24: o_data_a = 16'b1110110010100000;
            14'h3d25: o_data_a = 16'b1110001100001000;
            14'h3d26: o_data_a = 16'b0000000000110000;
            14'h3d27: o_data_a = 16'b1110110000010000;
            14'h3d28: o_data_a = 16'b0000000000000000;
            14'h3d29: o_data_a = 16'b1111110111101000;
            14'h3d2a: o_data_a = 16'b1110110010100000;
            14'h3d2b: o_data_a = 16'b1110001100001000;
            14'h3d2c: o_data_a = 16'b0000000000111100;
            14'h3d2d: o_data_a = 16'b1110110000010000;
            14'h3d2e: o_data_a = 16'b0000000000000000;
            14'h3d2f: o_data_a = 16'b1111110111101000;
            14'h3d30: o_data_a = 16'b1110110010100000;
            14'h3d31: o_data_a = 16'b1110001100001000;
            14'h3d32: o_data_a = 16'b0000000000110110;
            14'h3d33: o_data_a = 16'b1110110000010000;
            14'h3d34: o_data_a = 16'b0000000000000000;
            14'h3d35: o_data_a = 16'b1111110111101000;
            14'h3d36: o_data_a = 16'b1110110010100000;
            14'h3d37: o_data_a = 16'b1110001100001000;
            14'h3d38: o_data_a = 16'b0000000000110011;
            14'h3d39: o_data_a = 16'b1110110000010000;
            14'h3d3a: o_data_a = 16'b0000000000000000;
            14'h3d3b: o_data_a = 16'b1111110111101000;
            14'h3d3c: o_data_a = 16'b1110110010100000;
            14'h3d3d: o_data_a = 16'b1110001100001000;
            14'h3d3e: o_data_a = 16'b0000000000110011;
            14'h3d3f: o_data_a = 16'b1110110000010000;
            14'h3d40: o_data_a = 16'b0000000000000000;
            14'h3d41: o_data_a = 16'b1111110111101000;
            14'h3d42: o_data_a = 16'b1110110010100000;
            14'h3d43: o_data_a = 16'b1110001100001000;
            14'h3d44: o_data_a = 16'b0000000000110011;
            14'h3d45: o_data_a = 16'b1110110000010000;
            14'h3d46: o_data_a = 16'b0000000000000000;
            14'h3d47: o_data_a = 16'b1111110111101000;
            14'h3d48: o_data_a = 16'b1110110010100000;
            14'h3d49: o_data_a = 16'b1110001100001000;
            14'h3d4a: o_data_a = 16'b0000000000011110;
            14'h3d4b: o_data_a = 16'b1110110000010000;
            14'h3d4c: o_data_a = 16'b0000000000000000;
            14'h3d4d: o_data_a = 16'b1111110111101000;
            14'h3d4e: o_data_a = 16'b1110110010100000;
            14'h3d4f: o_data_a = 16'b1110001100001000;
            14'h3d50: o_data_a = 16'b0000000000000000;
            14'h3d51: o_data_a = 16'b1111110111001000;
            14'h3d52: o_data_a = 16'b1111110010100000;
            14'h3d53: o_data_a = 16'b1110101010001000;
            14'h3d54: o_data_a = 16'b0000000000000000;
            14'h3d55: o_data_a = 16'b1111110111001000;
            14'h3d56: o_data_a = 16'b1111110010100000;
            14'h3d57: o_data_a = 16'b1110101010001000;
            14'h3d58: o_data_a = 16'b0000000000001100;
            14'h3d59: o_data_a = 16'b1110110000010000;
            14'h3d5a: o_data_a = 16'b0000000000001101;
            14'h3d5b: o_data_a = 16'b1110001100001000;
            14'h3d5c: o_data_a = 16'b0100010110110011;
            14'h3d5d: o_data_a = 16'b1110110000010000;
            14'h3d5e: o_data_a = 16'b0000000000001110;
            14'h3d5f: o_data_a = 16'b1110001100001000;
            14'h3d60: o_data_a = 16'b0011110101100100;
            14'h3d61: o_data_a = 16'b1110110000010000;
            14'h3d62: o_data_a = 16'b0000000001011111;
            14'h3d63: o_data_a = 16'b1110101010000111;
            14'h3d64: o_data_a = 16'b0000000000000000;
            14'h3d65: o_data_a = 16'b1111110010101000;
            14'h3d66: o_data_a = 16'b1111110000010000;
            14'h3d67: o_data_a = 16'b0000000000000101;
            14'h3d68: o_data_a = 16'b1110001100001000;
            14'h3d69: o_data_a = 16'b0000000001100101;
            14'h3d6a: o_data_a = 16'b1110110000010000;
            14'h3d6b: o_data_a = 16'b0000000000000000;
            14'h3d6c: o_data_a = 16'b1111110111101000;
            14'h3d6d: o_data_a = 16'b1110110010100000;
            14'h3d6e: o_data_a = 16'b1110001100001000;
            14'h3d6f: o_data_a = 16'b0000000000000000;
            14'h3d70: o_data_a = 16'b1111110111001000;
            14'h3d71: o_data_a = 16'b1111110010100000;
            14'h3d72: o_data_a = 16'b1110101010001000;
            14'h3d73: o_data_a = 16'b0000000000000000;
            14'h3d74: o_data_a = 16'b1111110111001000;
            14'h3d75: o_data_a = 16'b1111110010100000;
            14'h3d76: o_data_a = 16'b1110101010001000;
            14'h3d77: o_data_a = 16'b0000000000000000;
            14'h3d78: o_data_a = 16'b1111110111001000;
            14'h3d79: o_data_a = 16'b1111110010100000;
            14'h3d7a: o_data_a = 16'b1110101010001000;
            14'h3d7b: o_data_a = 16'b0000000000011110;
            14'h3d7c: o_data_a = 16'b1110110000010000;
            14'h3d7d: o_data_a = 16'b0000000000000000;
            14'h3d7e: o_data_a = 16'b1111110111101000;
            14'h3d7f: o_data_a = 16'b1110110010100000;
            14'h3d80: o_data_a = 16'b1110001100001000;
            14'h3d81: o_data_a = 16'b0000000000110011;
            14'h3d82: o_data_a = 16'b1110110000010000;
            14'h3d83: o_data_a = 16'b0000000000000000;
            14'h3d84: o_data_a = 16'b1111110111101000;
            14'h3d85: o_data_a = 16'b1110110010100000;
            14'h3d86: o_data_a = 16'b1110001100001000;
            14'h3d87: o_data_a = 16'b0000000000111111;
            14'h3d88: o_data_a = 16'b1110110000010000;
            14'h3d89: o_data_a = 16'b0000000000000000;
            14'h3d8a: o_data_a = 16'b1111110111101000;
            14'h3d8b: o_data_a = 16'b1110110010100000;
            14'h3d8c: o_data_a = 16'b1110001100001000;
            14'h3d8d: o_data_a = 16'b0000000000000011;
            14'h3d8e: o_data_a = 16'b1110110000010000;
            14'h3d8f: o_data_a = 16'b0000000000000000;
            14'h3d90: o_data_a = 16'b1111110111101000;
            14'h3d91: o_data_a = 16'b1110110010100000;
            14'h3d92: o_data_a = 16'b1110001100001000;
            14'h3d93: o_data_a = 16'b0000000000110011;
            14'h3d94: o_data_a = 16'b1110110000010000;
            14'h3d95: o_data_a = 16'b0000000000000000;
            14'h3d96: o_data_a = 16'b1111110111101000;
            14'h3d97: o_data_a = 16'b1110110010100000;
            14'h3d98: o_data_a = 16'b1110001100001000;
            14'h3d99: o_data_a = 16'b0000000000011110;
            14'h3d9a: o_data_a = 16'b1110110000010000;
            14'h3d9b: o_data_a = 16'b0000000000000000;
            14'h3d9c: o_data_a = 16'b1111110111101000;
            14'h3d9d: o_data_a = 16'b1110110010100000;
            14'h3d9e: o_data_a = 16'b1110001100001000;
            14'h3d9f: o_data_a = 16'b0000000000000000;
            14'h3da0: o_data_a = 16'b1111110111001000;
            14'h3da1: o_data_a = 16'b1111110010100000;
            14'h3da2: o_data_a = 16'b1110101010001000;
            14'h3da3: o_data_a = 16'b0000000000000000;
            14'h3da4: o_data_a = 16'b1111110111001000;
            14'h3da5: o_data_a = 16'b1111110010100000;
            14'h3da6: o_data_a = 16'b1110101010001000;
            14'h3da7: o_data_a = 16'b0000000000001100;
            14'h3da8: o_data_a = 16'b1110110000010000;
            14'h3da9: o_data_a = 16'b0000000000001101;
            14'h3daa: o_data_a = 16'b1110001100001000;
            14'h3dab: o_data_a = 16'b0100010110110011;
            14'h3dac: o_data_a = 16'b1110110000010000;
            14'h3dad: o_data_a = 16'b0000000000001110;
            14'h3dae: o_data_a = 16'b1110001100001000;
            14'h3daf: o_data_a = 16'b0011110110110011;
            14'h3db0: o_data_a = 16'b1110110000010000;
            14'h3db1: o_data_a = 16'b0000000001011111;
            14'h3db2: o_data_a = 16'b1110101010000111;
            14'h3db3: o_data_a = 16'b0000000000000000;
            14'h3db4: o_data_a = 16'b1111110010101000;
            14'h3db5: o_data_a = 16'b1111110000010000;
            14'h3db6: o_data_a = 16'b0000000000000101;
            14'h3db7: o_data_a = 16'b1110001100001000;
            14'h3db8: o_data_a = 16'b0000000001100110;
            14'h3db9: o_data_a = 16'b1110110000010000;
            14'h3dba: o_data_a = 16'b0000000000000000;
            14'h3dbb: o_data_a = 16'b1111110111101000;
            14'h3dbc: o_data_a = 16'b1110110010100000;
            14'h3dbd: o_data_a = 16'b1110001100001000;
            14'h3dbe: o_data_a = 16'b0000000000011100;
            14'h3dbf: o_data_a = 16'b1110110000010000;
            14'h3dc0: o_data_a = 16'b0000000000000000;
            14'h3dc1: o_data_a = 16'b1111110111101000;
            14'h3dc2: o_data_a = 16'b1110110010100000;
            14'h3dc3: o_data_a = 16'b1110001100001000;
            14'h3dc4: o_data_a = 16'b0000000000110110;
            14'h3dc5: o_data_a = 16'b1110110000010000;
            14'h3dc6: o_data_a = 16'b0000000000000000;
            14'h3dc7: o_data_a = 16'b1111110111101000;
            14'h3dc8: o_data_a = 16'b1110110010100000;
            14'h3dc9: o_data_a = 16'b1110001100001000;
            14'h3dca: o_data_a = 16'b0000000000100110;
            14'h3dcb: o_data_a = 16'b1110110000010000;
            14'h3dcc: o_data_a = 16'b0000000000000000;
            14'h3dcd: o_data_a = 16'b1111110111101000;
            14'h3dce: o_data_a = 16'b1110110010100000;
            14'h3dcf: o_data_a = 16'b1110001100001000;
            14'h3dd0: o_data_a = 16'b0000000000000110;
            14'h3dd1: o_data_a = 16'b1110110000010000;
            14'h3dd2: o_data_a = 16'b0000000000000000;
            14'h3dd3: o_data_a = 16'b1111110111101000;
            14'h3dd4: o_data_a = 16'b1110110010100000;
            14'h3dd5: o_data_a = 16'b1110001100001000;
            14'h3dd6: o_data_a = 16'b0000000000001111;
            14'h3dd7: o_data_a = 16'b1110110000010000;
            14'h3dd8: o_data_a = 16'b0000000000000000;
            14'h3dd9: o_data_a = 16'b1111110111101000;
            14'h3dda: o_data_a = 16'b1110110010100000;
            14'h3ddb: o_data_a = 16'b1110001100001000;
            14'h3ddc: o_data_a = 16'b0000000000000110;
            14'h3ddd: o_data_a = 16'b1110110000010000;
            14'h3dde: o_data_a = 16'b0000000000000000;
            14'h3ddf: o_data_a = 16'b1111110111101000;
            14'h3de0: o_data_a = 16'b1110110010100000;
            14'h3de1: o_data_a = 16'b1110001100001000;
            14'h3de2: o_data_a = 16'b0000000000000110;
            14'h3de3: o_data_a = 16'b1110110000010000;
            14'h3de4: o_data_a = 16'b0000000000000000;
            14'h3de5: o_data_a = 16'b1111110111101000;
            14'h3de6: o_data_a = 16'b1110110010100000;
            14'h3de7: o_data_a = 16'b1110001100001000;
            14'h3de8: o_data_a = 16'b0000000000000110;
            14'h3de9: o_data_a = 16'b1110110000010000;
            14'h3dea: o_data_a = 16'b0000000000000000;
            14'h3deb: o_data_a = 16'b1111110111101000;
            14'h3dec: o_data_a = 16'b1110110010100000;
            14'h3ded: o_data_a = 16'b1110001100001000;
            14'h3dee: o_data_a = 16'b0000000000001111;
            14'h3def: o_data_a = 16'b1110110000010000;
            14'h3df0: o_data_a = 16'b0000000000000000;
            14'h3df1: o_data_a = 16'b1111110111101000;
            14'h3df2: o_data_a = 16'b1110110010100000;
            14'h3df3: o_data_a = 16'b1110001100001000;
            14'h3df4: o_data_a = 16'b0000000000000000;
            14'h3df5: o_data_a = 16'b1111110111001000;
            14'h3df6: o_data_a = 16'b1111110010100000;
            14'h3df7: o_data_a = 16'b1110101010001000;
            14'h3df8: o_data_a = 16'b0000000000000000;
            14'h3df9: o_data_a = 16'b1111110111001000;
            14'h3dfa: o_data_a = 16'b1111110010100000;
            14'h3dfb: o_data_a = 16'b1110101010001000;
            14'h3dfc: o_data_a = 16'b0000000000001100;
            14'h3dfd: o_data_a = 16'b1110110000010000;
            14'h3dfe: o_data_a = 16'b0000000000001101;
            14'h3dff: o_data_a = 16'b1110001100001000;
            14'h3e00: o_data_a = 16'b0100010110110011;
            14'h3e01: o_data_a = 16'b1110110000010000;
            14'h3e02: o_data_a = 16'b0000000000001110;
            14'h3e03: o_data_a = 16'b1110001100001000;
            14'h3e04: o_data_a = 16'b0011111000001000;
            14'h3e05: o_data_a = 16'b1110110000010000;
            14'h3e06: o_data_a = 16'b0000000001011111;
            14'h3e07: o_data_a = 16'b1110101010000111;
            14'h3e08: o_data_a = 16'b0000000000000000;
            14'h3e09: o_data_a = 16'b1111110010101000;
            14'h3e0a: o_data_a = 16'b1111110000010000;
            14'h3e0b: o_data_a = 16'b0000000000000101;
            14'h3e0c: o_data_a = 16'b1110001100001000;
            14'h3e0d: o_data_a = 16'b0000000001100111;
            14'h3e0e: o_data_a = 16'b1110110000010000;
            14'h3e0f: o_data_a = 16'b0000000000000000;
            14'h3e10: o_data_a = 16'b1111110111101000;
            14'h3e11: o_data_a = 16'b1110110010100000;
            14'h3e12: o_data_a = 16'b1110001100001000;
            14'h3e13: o_data_a = 16'b0000000000000000;
            14'h3e14: o_data_a = 16'b1111110111001000;
            14'h3e15: o_data_a = 16'b1111110010100000;
            14'h3e16: o_data_a = 16'b1110101010001000;
            14'h3e17: o_data_a = 16'b0000000000000000;
            14'h3e18: o_data_a = 16'b1111110111001000;
            14'h3e19: o_data_a = 16'b1111110010100000;
            14'h3e1a: o_data_a = 16'b1110101010001000;
            14'h3e1b: o_data_a = 16'b0000000000011110;
            14'h3e1c: o_data_a = 16'b1110110000010000;
            14'h3e1d: o_data_a = 16'b0000000000000000;
            14'h3e1e: o_data_a = 16'b1111110111101000;
            14'h3e1f: o_data_a = 16'b1110110010100000;
            14'h3e20: o_data_a = 16'b1110001100001000;
            14'h3e21: o_data_a = 16'b0000000000110011;
            14'h3e22: o_data_a = 16'b1110110000010000;
            14'h3e23: o_data_a = 16'b0000000000000000;
            14'h3e24: o_data_a = 16'b1111110111101000;
            14'h3e25: o_data_a = 16'b1110110010100000;
            14'h3e26: o_data_a = 16'b1110001100001000;
            14'h3e27: o_data_a = 16'b0000000000110011;
            14'h3e28: o_data_a = 16'b1110110000010000;
            14'h3e29: o_data_a = 16'b0000000000000000;
            14'h3e2a: o_data_a = 16'b1111110111101000;
            14'h3e2b: o_data_a = 16'b1110110010100000;
            14'h3e2c: o_data_a = 16'b1110001100001000;
            14'h3e2d: o_data_a = 16'b0000000000110011;
            14'h3e2e: o_data_a = 16'b1110110000010000;
            14'h3e2f: o_data_a = 16'b0000000000000000;
            14'h3e30: o_data_a = 16'b1111110111101000;
            14'h3e31: o_data_a = 16'b1110110010100000;
            14'h3e32: o_data_a = 16'b1110001100001000;
            14'h3e33: o_data_a = 16'b0000000000111110;
            14'h3e34: o_data_a = 16'b1110110000010000;
            14'h3e35: o_data_a = 16'b0000000000000000;
            14'h3e36: o_data_a = 16'b1111110111101000;
            14'h3e37: o_data_a = 16'b1110110010100000;
            14'h3e38: o_data_a = 16'b1110001100001000;
            14'h3e39: o_data_a = 16'b0000000000110000;
            14'h3e3a: o_data_a = 16'b1110110000010000;
            14'h3e3b: o_data_a = 16'b0000000000000000;
            14'h3e3c: o_data_a = 16'b1111110111101000;
            14'h3e3d: o_data_a = 16'b1110110010100000;
            14'h3e3e: o_data_a = 16'b1110001100001000;
            14'h3e3f: o_data_a = 16'b0000000000110011;
            14'h3e40: o_data_a = 16'b1110110000010000;
            14'h3e41: o_data_a = 16'b0000000000000000;
            14'h3e42: o_data_a = 16'b1111110111101000;
            14'h3e43: o_data_a = 16'b1110110010100000;
            14'h3e44: o_data_a = 16'b1110001100001000;
            14'h3e45: o_data_a = 16'b0000000000011110;
            14'h3e46: o_data_a = 16'b1110110000010000;
            14'h3e47: o_data_a = 16'b0000000000000000;
            14'h3e48: o_data_a = 16'b1111110111101000;
            14'h3e49: o_data_a = 16'b1110110010100000;
            14'h3e4a: o_data_a = 16'b1110001100001000;
            14'h3e4b: o_data_a = 16'b0000000000000000;
            14'h3e4c: o_data_a = 16'b1111110111001000;
            14'h3e4d: o_data_a = 16'b1111110010100000;
            14'h3e4e: o_data_a = 16'b1110101010001000;
            14'h3e4f: o_data_a = 16'b0000000000001100;
            14'h3e50: o_data_a = 16'b1110110000010000;
            14'h3e51: o_data_a = 16'b0000000000001101;
            14'h3e52: o_data_a = 16'b1110001100001000;
            14'h3e53: o_data_a = 16'b0100010110110011;
            14'h3e54: o_data_a = 16'b1110110000010000;
            14'h3e55: o_data_a = 16'b0000000000001110;
            14'h3e56: o_data_a = 16'b1110001100001000;
            14'h3e57: o_data_a = 16'b0011111001011011;
            14'h3e58: o_data_a = 16'b1110110000010000;
            14'h3e59: o_data_a = 16'b0000000001011111;
            14'h3e5a: o_data_a = 16'b1110101010000111;
            14'h3e5b: o_data_a = 16'b0000000000000000;
            14'h3e5c: o_data_a = 16'b1111110010101000;
            14'h3e5d: o_data_a = 16'b1111110000010000;
            14'h3e5e: o_data_a = 16'b0000000000000101;
            14'h3e5f: o_data_a = 16'b1110001100001000;
            14'h3e60: o_data_a = 16'b0000000001101000;
            14'h3e61: o_data_a = 16'b1110110000010000;
            14'h3e62: o_data_a = 16'b0000000000000000;
            14'h3e63: o_data_a = 16'b1111110111101000;
            14'h3e64: o_data_a = 16'b1110110010100000;
            14'h3e65: o_data_a = 16'b1110001100001000;
            14'h3e66: o_data_a = 16'b0000000000000011;
            14'h3e67: o_data_a = 16'b1110110000010000;
            14'h3e68: o_data_a = 16'b0000000000000000;
            14'h3e69: o_data_a = 16'b1111110111101000;
            14'h3e6a: o_data_a = 16'b1110110010100000;
            14'h3e6b: o_data_a = 16'b1110001100001000;
            14'h3e6c: o_data_a = 16'b0000000000000011;
            14'h3e6d: o_data_a = 16'b1110110000010000;
            14'h3e6e: o_data_a = 16'b0000000000000000;
            14'h3e6f: o_data_a = 16'b1111110111101000;
            14'h3e70: o_data_a = 16'b1110110010100000;
            14'h3e71: o_data_a = 16'b1110001100001000;
            14'h3e72: o_data_a = 16'b0000000000000011;
            14'h3e73: o_data_a = 16'b1110110000010000;
            14'h3e74: o_data_a = 16'b0000000000000000;
            14'h3e75: o_data_a = 16'b1111110111101000;
            14'h3e76: o_data_a = 16'b1110110010100000;
            14'h3e77: o_data_a = 16'b1110001100001000;
            14'h3e78: o_data_a = 16'b0000000000011011;
            14'h3e79: o_data_a = 16'b1110110000010000;
            14'h3e7a: o_data_a = 16'b0000000000000000;
            14'h3e7b: o_data_a = 16'b1111110111101000;
            14'h3e7c: o_data_a = 16'b1110110010100000;
            14'h3e7d: o_data_a = 16'b1110001100001000;
            14'h3e7e: o_data_a = 16'b0000000000110111;
            14'h3e7f: o_data_a = 16'b1110110000010000;
            14'h3e80: o_data_a = 16'b0000000000000000;
            14'h3e81: o_data_a = 16'b1111110111101000;
            14'h3e82: o_data_a = 16'b1110110010100000;
            14'h3e83: o_data_a = 16'b1110001100001000;
            14'h3e84: o_data_a = 16'b0000000000110011;
            14'h3e85: o_data_a = 16'b1110110000010000;
            14'h3e86: o_data_a = 16'b0000000000000000;
            14'h3e87: o_data_a = 16'b1111110111101000;
            14'h3e88: o_data_a = 16'b1110110010100000;
            14'h3e89: o_data_a = 16'b1110001100001000;
            14'h3e8a: o_data_a = 16'b0000000000110011;
            14'h3e8b: o_data_a = 16'b1110110000010000;
            14'h3e8c: o_data_a = 16'b0000000000000000;
            14'h3e8d: o_data_a = 16'b1111110111101000;
            14'h3e8e: o_data_a = 16'b1110110010100000;
            14'h3e8f: o_data_a = 16'b1110001100001000;
            14'h3e90: o_data_a = 16'b0000000000110011;
            14'h3e91: o_data_a = 16'b1110110000010000;
            14'h3e92: o_data_a = 16'b0000000000000000;
            14'h3e93: o_data_a = 16'b1111110111101000;
            14'h3e94: o_data_a = 16'b1110110010100000;
            14'h3e95: o_data_a = 16'b1110001100001000;
            14'h3e96: o_data_a = 16'b0000000000110011;
            14'h3e97: o_data_a = 16'b1110110000010000;
            14'h3e98: o_data_a = 16'b0000000000000000;
            14'h3e99: o_data_a = 16'b1111110111101000;
            14'h3e9a: o_data_a = 16'b1110110010100000;
            14'h3e9b: o_data_a = 16'b1110001100001000;
            14'h3e9c: o_data_a = 16'b0000000000000000;
            14'h3e9d: o_data_a = 16'b1111110111001000;
            14'h3e9e: o_data_a = 16'b1111110010100000;
            14'h3e9f: o_data_a = 16'b1110101010001000;
            14'h3ea0: o_data_a = 16'b0000000000000000;
            14'h3ea1: o_data_a = 16'b1111110111001000;
            14'h3ea2: o_data_a = 16'b1111110010100000;
            14'h3ea3: o_data_a = 16'b1110101010001000;
            14'h3ea4: o_data_a = 16'b0000000000001100;
            14'h3ea5: o_data_a = 16'b1110110000010000;
            14'h3ea6: o_data_a = 16'b0000000000001101;
            14'h3ea7: o_data_a = 16'b1110001100001000;
            14'h3ea8: o_data_a = 16'b0100010110110011;
            14'h3ea9: o_data_a = 16'b1110110000010000;
            14'h3eaa: o_data_a = 16'b0000000000001110;
            14'h3eab: o_data_a = 16'b1110001100001000;
            14'h3eac: o_data_a = 16'b0011111010110000;
            14'h3ead: o_data_a = 16'b1110110000010000;
            14'h3eae: o_data_a = 16'b0000000001011111;
            14'h3eaf: o_data_a = 16'b1110101010000111;
            14'h3eb0: o_data_a = 16'b0000000000000000;
            14'h3eb1: o_data_a = 16'b1111110010101000;
            14'h3eb2: o_data_a = 16'b1111110000010000;
            14'h3eb3: o_data_a = 16'b0000000000000101;
            14'h3eb4: o_data_a = 16'b1110001100001000;
            14'h3eb5: o_data_a = 16'b0000000001101001;
            14'h3eb6: o_data_a = 16'b1110110000010000;
            14'h3eb7: o_data_a = 16'b0000000000000000;
            14'h3eb8: o_data_a = 16'b1111110111101000;
            14'h3eb9: o_data_a = 16'b1110110010100000;
            14'h3eba: o_data_a = 16'b1110001100001000;
            14'h3ebb: o_data_a = 16'b0000000000001100;
            14'h3ebc: o_data_a = 16'b1110110000010000;
            14'h3ebd: o_data_a = 16'b0000000000000000;
            14'h3ebe: o_data_a = 16'b1111110111101000;
            14'h3ebf: o_data_a = 16'b1110110010100000;
            14'h3ec0: o_data_a = 16'b1110001100001000;
            14'h3ec1: o_data_a = 16'b0000000000001100;
            14'h3ec2: o_data_a = 16'b1110110000010000;
            14'h3ec3: o_data_a = 16'b0000000000000000;
            14'h3ec4: o_data_a = 16'b1111110111101000;
            14'h3ec5: o_data_a = 16'b1110110010100000;
            14'h3ec6: o_data_a = 16'b1110001100001000;
            14'h3ec7: o_data_a = 16'b0000000000000000;
            14'h3ec8: o_data_a = 16'b1111110111001000;
            14'h3ec9: o_data_a = 16'b1111110010100000;
            14'h3eca: o_data_a = 16'b1110101010001000;
            14'h3ecb: o_data_a = 16'b0000000000001110;
            14'h3ecc: o_data_a = 16'b1110110000010000;
            14'h3ecd: o_data_a = 16'b0000000000000000;
            14'h3ece: o_data_a = 16'b1111110111101000;
            14'h3ecf: o_data_a = 16'b1110110010100000;
            14'h3ed0: o_data_a = 16'b1110001100001000;
            14'h3ed1: o_data_a = 16'b0000000000001100;
            14'h3ed2: o_data_a = 16'b1110110000010000;
            14'h3ed3: o_data_a = 16'b0000000000000000;
            14'h3ed4: o_data_a = 16'b1111110111101000;
            14'h3ed5: o_data_a = 16'b1110110010100000;
            14'h3ed6: o_data_a = 16'b1110001100001000;
            14'h3ed7: o_data_a = 16'b0000000000001100;
            14'h3ed8: o_data_a = 16'b1110110000010000;
            14'h3ed9: o_data_a = 16'b0000000000000000;
            14'h3eda: o_data_a = 16'b1111110111101000;
            14'h3edb: o_data_a = 16'b1110110010100000;
            14'h3edc: o_data_a = 16'b1110001100001000;
            14'h3edd: o_data_a = 16'b0000000000001100;
            14'h3ede: o_data_a = 16'b1110110000010000;
            14'h3edf: o_data_a = 16'b0000000000000000;
            14'h3ee0: o_data_a = 16'b1111110111101000;
            14'h3ee1: o_data_a = 16'b1110110010100000;
            14'h3ee2: o_data_a = 16'b1110001100001000;
            14'h3ee3: o_data_a = 16'b0000000000001100;
            14'h3ee4: o_data_a = 16'b1110110000010000;
            14'h3ee5: o_data_a = 16'b0000000000000000;
            14'h3ee6: o_data_a = 16'b1111110111101000;
            14'h3ee7: o_data_a = 16'b1110110010100000;
            14'h3ee8: o_data_a = 16'b1110001100001000;
            14'h3ee9: o_data_a = 16'b0000000000011110;
            14'h3eea: o_data_a = 16'b1110110000010000;
            14'h3eeb: o_data_a = 16'b0000000000000000;
            14'h3eec: o_data_a = 16'b1111110111101000;
            14'h3eed: o_data_a = 16'b1110110010100000;
            14'h3eee: o_data_a = 16'b1110001100001000;
            14'h3eef: o_data_a = 16'b0000000000000000;
            14'h3ef0: o_data_a = 16'b1111110111001000;
            14'h3ef1: o_data_a = 16'b1111110010100000;
            14'h3ef2: o_data_a = 16'b1110101010001000;
            14'h3ef3: o_data_a = 16'b0000000000000000;
            14'h3ef4: o_data_a = 16'b1111110111001000;
            14'h3ef5: o_data_a = 16'b1111110010100000;
            14'h3ef6: o_data_a = 16'b1110101010001000;
            14'h3ef7: o_data_a = 16'b0000000000001100;
            14'h3ef8: o_data_a = 16'b1110110000010000;
            14'h3ef9: o_data_a = 16'b0000000000001101;
            14'h3efa: o_data_a = 16'b1110001100001000;
            14'h3efb: o_data_a = 16'b0100010110110011;
            14'h3efc: o_data_a = 16'b1110110000010000;
            14'h3efd: o_data_a = 16'b0000000000001110;
            14'h3efe: o_data_a = 16'b1110001100001000;
            14'h3eff: o_data_a = 16'b0011111100000011;
            14'h3f00: o_data_a = 16'b1110110000010000;
            14'h3f01: o_data_a = 16'b0000000001011111;
            14'h3f02: o_data_a = 16'b1110101010000111;
            14'h3f03: o_data_a = 16'b0000000000000000;
            14'h3f04: o_data_a = 16'b1111110010101000;
            14'h3f05: o_data_a = 16'b1111110000010000;
            14'h3f06: o_data_a = 16'b0000000000000101;
            14'h3f07: o_data_a = 16'b1110001100001000;
            14'h3f08: o_data_a = 16'b0000000001101010;
            14'h3f09: o_data_a = 16'b1110110000010000;
            14'h3f0a: o_data_a = 16'b0000000000000000;
            14'h3f0b: o_data_a = 16'b1111110111101000;
            14'h3f0c: o_data_a = 16'b1110110010100000;
            14'h3f0d: o_data_a = 16'b1110001100001000;
            14'h3f0e: o_data_a = 16'b0000000000110000;
            14'h3f0f: o_data_a = 16'b1110110000010000;
            14'h3f10: o_data_a = 16'b0000000000000000;
            14'h3f11: o_data_a = 16'b1111110111101000;
            14'h3f12: o_data_a = 16'b1110110010100000;
            14'h3f13: o_data_a = 16'b1110001100001000;
            14'h3f14: o_data_a = 16'b0000000000110000;
            14'h3f15: o_data_a = 16'b1110110000010000;
            14'h3f16: o_data_a = 16'b0000000000000000;
            14'h3f17: o_data_a = 16'b1111110111101000;
            14'h3f18: o_data_a = 16'b1110110010100000;
            14'h3f19: o_data_a = 16'b1110001100001000;
            14'h3f1a: o_data_a = 16'b0000000000000000;
            14'h3f1b: o_data_a = 16'b1111110111001000;
            14'h3f1c: o_data_a = 16'b1111110010100000;
            14'h3f1d: o_data_a = 16'b1110101010001000;
            14'h3f1e: o_data_a = 16'b0000000000111000;
            14'h3f1f: o_data_a = 16'b1110110000010000;
            14'h3f20: o_data_a = 16'b0000000000000000;
            14'h3f21: o_data_a = 16'b1111110111101000;
            14'h3f22: o_data_a = 16'b1110110010100000;
            14'h3f23: o_data_a = 16'b1110001100001000;
            14'h3f24: o_data_a = 16'b0000000000110000;
            14'h3f25: o_data_a = 16'b1110110000010000;
            14'h3f26: o_data_a = 16'b0000000000000000;
            14'h3f27: o_data_a = 16'b1111110111101000;
            14'h3f28: o_data_a = 16'b1110110010100000;
            14'h3f29: o_data_a = 16'b1110001100001000;
            14'h3f2a: o_data_a = 16'b0000000000110000;
            14'h3f2b: o_data_a = 16'b1110110000010000;
            14'h3f2c: o_data_a = 16'b0000000000000000;
            14'h3f2d: o_data_a = 16'b1111110111101000;
            14'h3f2e: o_data_a = 16'b1110110010100000;
            14'h3f2f: o_data_a = 16'b1110001100001000;
            14'h3f30: o_data_a = 16'b0000000000110000;
            14'h3f31: o_data_a = 16'b1110110000010000;
            14'h3f32: o_data_a = 16'b0000000000000000;
            14'h3f33: o_data_a = 16'b1111110111101000;
            14'h3f34: o_data_a = 16'b1110110010100000;
            14'h3f35: o_data_a = 16'b1110001100001000;
            14'h3f36: o_data_a = 16'b0000000000110000;
            14'h3f37: o_data_a = 16'b1110110000010000;
            14'h3f38: o_data_a = 16'b0000000000000000;
            14'h3f39: o_data_a = 16'b1111110111101000;
            14'h3f3a: o_data_a = 16'b1110110010100000;
            14'h3f3b: o_data_a = 16'b1110001100001000;
            14'h3f3c: o_data_a = 16'b0000000000110011;
            14'h3f3d: o_data_a = 16'b1110110000010000;
            14'h3f3e: o_data_a = 16'b0000000000000000;
            14'h3f3f: o_data_a = 16'b1111110111101000;
            14'h3f40: o_data_a = 16'b1110110010100000;
            14'h3f41: o_data_a = 16'b1110001100001000;
            14'h3f42: o_data_a = 16'b0000000000011110;
            14'h3f43: o_data_a = 16'b1110110000010000;
            14'h3f44: o_data_a = 16'b0000000000000000;
            14'h3f45: o_data_a = 16'b1111110111101000;
            14'h3f46: o_data_a = 16'b1110110010100000;
            14'h3f47: o_data_a = 16'b1110001100001000;
            14'h3f48: o_data_a = 16'b0000000000000000;
            14'h3f49: o_data_a = 16'b1111110111001000;
            14'h3f4a: o_data_a = 16'b1111110010100000;
            14'h3f4b: o_data_a = 16'b1110101010001000;
            14'h3f4c: o_data_a = 16'b0000000000001100;
            14'h3f4d: o_data_a = 16'b1110110000010000;
            14'h3f4e: o_data_a = 16'b0000000000001101;
            14'h3f4f: o_data_a = 16'b1110001100001000;
            14'h3f50: o_data_a = 16'b0100010110110011;
            14'h3f51: o_data_a = 16'b1110110000010000;
            14'h3f52: o_data_a = 16'b0000000000001110;
            14'h3f53: o_data_a = 16'b1110001100001000;
            14'h3f54: o_data_a = 16'b0011111101011000;
            14'h3f55: o_data_a = 16'b1110110000010000;
            14'h3f56: o_data_a = 16'b0000000001011111;
            14'h3f57: o_data_a = 16'b1110101010000111;
            14'h3f58: o_data_a = 16'b0000000000000000;
            14'h3f59: o_data_a = 16'b1111110010101000;
            14'h3f5a: o_data_a = 16'b1111110000010000;
            14'h3f5b: o_data_a = 16'b0000000000000101;
            14'h3f5c: o_data_a = 16'b1110001100001000;
            14'h3f5d: o_data_a = 16'b0000000001101011;
            14'h3f5e: o_data_a = 16'b1110110000010000;
            14'h3f5f: o_data_a = 16'b0000000000000000;
            14'h3f60: o_data_a = 16'b1111110111101000;
            14'h3f61: o_data_a = 16'b1110110010100000;
            14'h3f62: o_data_a = 16'b1110001100001000;
            14'h3f63: o_data_a = 16'b0000000000000011;
            14'h3f64: o_data_a = 16'b1110110000010000;
            14'h3f65: o_data_a = 16'b0000000000000000;
            14'h3f66: o_data_a = 16'b1111110111101000;
            14'h3f67: o_data_a = 16'b1110110010100000;
            14'h3f68: o_data_a = 16'b1110001100001000;
            14'h3f69: o_data_a = 16'b0000000000000011;
            14'h3f6a: o_data_a = 16'b1110110000010000;
            14'h3f6b: o_data_a = 16'b0000000000000000;
            14'h3f6c: o_data_a = 16'b1111110111101000;
            14'h3f6d: o_data_a = 16'b1110110010100000;
            14'h3f6e: o_data_a = 16'b1110001100001000;
            14'h3f6f: o_data_a = 16'b0000000000000011;
            14'h3f70: o_data_a = 16'b1110110000010000;
            14'h3f71: o_data_a = 16'b0000000000000000;
            14'h3f72: o_data_a = 16'b1111110111101000;
            14'h3f73: o_data_a = 16'b1110110010100000;
            14'h3f74: o_data_a = 16'b1110001100001000;
            14'h3f75: o_data_a = 16'b0000000000110011;
            14'h3f76: o_data_a = 16'b1110110000010000;
            14'h3f77: o_data_a = 16'b0000000000000000;
            14'h3f78: o_data_a = 16'b1111110111101000;
            14'h3f79: o_data_a = 16'b1110110010100000;
            14'h3f7a: o_data_a = 16'b1110001100001000;
            14'h3f7b: o_data_a = 16'b0000000000011011;
            14'h3f7c: o_data_a = 16'b1110110000010000;
            14'h3f7d: o_data_a = 16'b0000000000000000;
            14'h3f7e: o_data_a = 16'b1111110111101000;
            14'h3f7f: o_data_a = 16'b1110110010100000;
            14'h3f80: o_data_a = 16'b1110001100001000;
            14'h3f81: o_data_a = 16'b0000000000001111;
            14'h3f82: o_data_a = 16'b1110110000010000;
            14'h3f83: o_data_a = 16'b0000000000000000;
            14'h3f84: o_data_a = 16'b1111110111101000;
            14'h3f85: o_data_a = 16'b1110110010100000;
            14'h3f86: o_data_a = 16'b1110001100001000;
            14'h3f87: o_data_a = 16'b0000000000001111;
            14'h3f88: o_data_a = 16'b1110110000010000;
            14'h3f89: o_data_a = 16'b0000000000000000;
            14'h3f8a: o_data_a = 16'b1111110111101000;
            14'h3f8b: o_data_a = 16'b1110110010100000;
            14'h3f8c: o_data_a = 16'b1110001100001000;
            14'h3f8d: o_data_a = 16'b0000000000011011;
            14'h3f8e: o_data_a = 16'b1110110000010000;
            14'h3f8f: o_data_a = 16'b0000000000000000;
            14'h3f90: o_data_a = 16'b1111110111101000;
            14'h3f91: o_data_a = 16'b1110110010100000;
            14'h3f92: o_data_a = 16'b1110001100001000;
            14'h3f93: o_data_a = 16'b0000000000110011;
            14'h3f94: o_data_a = 16'b1110110000010000;
            14'h3f95: o_data_a = 16'b0000000000000000;
            14'h3f96: o_data_a = 16'b1111110111101000;
            14'h3f97: o_data_a = 16'b1110110010100000;
            14'h3f98: o_data_a = 16'b1110001100001000;
            14'h3f99: o_data_a = 16'b0000000000000000;
            14'h3f9a: o_data_a = 16'b1111110111001000;
            14'h3f9b: o_data_a = 16'b1111110010100000;
            14'h3f9c: o_data_a = 16'b1110101010001000;
            14'h3f9d: o_data_a = 16'b0000000000000000;
            14'h3f9e: o_data_a = 16'b1111110111001000;
            14'h3f9f: o_data_a = 16'b1111110010100000;
            14'h3fa0: o_data_a = 16'b1110101010001000;
            14'h3fa1: o_data_a = 16'b0000000000001100;
            14'h3fa2: o_data_a = 16'b1110110000010000;
            14'h3fa3: o_data_a = 16'b0000000000001101;
            14'h3fa4: o_data_a = 16'b1110001100001000;
            14'h3fa5: o_data_a = 16'b0100010110110011;
            14'h3fa6: o_data_a = 16'b1110110000010000;
            14'h3fa7: o_data_a = 16'b0000000000001110;
            14'h3fa8: o_data_a = 16'b1110001100001000;
            14'h3fa9: o_data_a = 16'b0011111110101101;
            14'h3faa: o_data_a = 16'b1110110000010000;
            14'h3fab: o_data_a = 16'b0000000001011111;
            14'h3fac: o_data_a = 16'b1110101010000111;
            14'h3fad: o_data_a = 16'b0000000000000000;
            14'h3fae: o_data_a = 16'b1111110010101000;
            14'h3faf: o_data_a = 16'b1111110000010000;
            14'h3fb0: o_data_a = 16'b0000000000000101;
            14'h3fb1: o_data_a = 16'b1110001100001000;
            14'h3fb2: o_data_a = 16'b0000000001101100;
            14'h3fb3: o_data_a = 16'b1110110000010000;
            14'h3fb4: o_data_a = 16'b0000000000000000;
            14'h3fb5: o_data_a = 16'b1111110111101000;
            14'h3fb6: o_data_a = 16'b1110110010100000;
            14'h3fb7: o_data_a = 16'b1110001100001000;
            14'h3fb8: o_data_a = 16'b0000000000001110;
            14'h3fb9: o_data_a = 16'b1110110000010000;
            14'h3fba: o_data_a = 16'b0000000000000000;
            14'h3fbb: o_data_a = 16'b1111110111101000;
            14'h3fbc: o_data_a = 16'b1110110010100000;
            14'h3fbd: o_data_a = 16'b1110001100001000;
            14'h3fbe: o_data_a = 16'b0000000000001100;
            14'h3fbf: o_data_a = 16'b1110110000010000;
            14'h3fc0: o_data_a = 16'b0000000000000000;
            14'h3fc1: o_data_a = 16'b1111110111101000;
            14'h3fc2: o_data_a = 16'b1110110010100000;
            14'h3fc3: o_data_a = 16'b1110001100001000;
            14'h3fc4: o_data_a = 16'b0000000000001100;
            14'h3fc5: o_data_a = 16'b1110110000010000;
            14'h3fc6: o_data_a = 16'b0000000000000000;
            14'h3fc7: o_data_a = 16'b1111110111101000;
            14'h3fc8: o_data_a = 16'b1110110010100000;
            14'h3fc9: o_data_a = 16'b1110001100001000;
            14'h3fca: o_data_a = 16'b0000000000001100;
            14'h3fcb: o_data_a = 16'b1110110000010000;
            14'h3fcc: o_data_a = 16'b0000000000000000;
            14'h3fcd: o_data_a = 16'b1111110111101000;
            14'h3fce: o_data_a = 16'b1110110010100000;
            14'h3fcf: o_data_a = 16'b1110001100001000;
            14'h3fd0: o_data_a = 16'b0000000000001100;
            14'h3fd1: o_data_a = 16'b1110110000010000;
            14'h3fd2: o_data_a = 16'b0000000000000000;
            14'h3fd3: o_data_a = 16'b1111110111101000;
            14'h3fd4: o_data_a = 16'b1110110010100000;
            14'h3fd5: o_data_a = 16'b1110001100001000;
            14'h3fd6: o_data_a = 16'b0000000000001100;
            14'h3fd7: o_data_a = 16'b1110110000010000;
            14'h3fd8: o_data_a = 16'b0000000000000000;
            14'h3fd9: o_data_a = 16'b1111110111101000;
            14'h3fda: o_data_a = 16'b1110110010100000;
            14'h3fdb: o_data_a = 16'b1110001100001000;
            14'h3fdc: o_data_a = 16'b0000000000001100;
            14'h3fdd: o_data_a = 16'b1110110000010000;
            14'h3fde: o_data_a = 16'b0000000000000000;
            14'h3fdf: o_data_a = 16'b1111110111101000;
            14'h3fe0: o_data_a = 16'b1110110010100000;
            14'h3fe1: o_data_a = 16'b1110001100001000;
            14'h3fe2: o_data_a = 16'b0000000000001100;
            14'h3fe3: o_data_a = 16'b1110110000010000;
            14'h3fe4: o_data_a = 16'b0000000000000000;
            14'h3fe5: o_data_a = 16'b1111110111101000;
            14'h3fe6: o_data_a = 16'b1110110010100000;
            14'h3fe7: o_data_a = 16'b1110001100001000;
            14'h3fe8: o_data_a = 16'b0000000000011110;
            14'h3fe9: o_data_a = 16'b1110110000010000;
            14'h3fea: o_data_a = 16'b0000000000000000;
            14'h3feb: o_data_a = 16'b1111110111101000;
            14'h3fec: o_data_a = 16'b1110110010100000;
            14'h3fed: o_data_a = 16'b1110001100001000;
            14'h3fee: o_data_a = 16'b0000000000000000;
            14'h3fef: o_data_a = 16'b1111110111001000;
            14'h3ff0: o_data_a = 16'b1111110010100000;
            14'h3ff1: o_data_a = 16'b1110101010001000;
            14'h3ff2: o_data_a = 16'b0000000000000000;
            14'h3ff3: o_data_a = 16'b1111110111001000;
            14'h3ff4: o_data_a = 16'b1111110010100000;
            14'h3ff5: o_data_a = 16'b1110101010001000;
            14'h3ff6: o_data_a = 16'b0000000000001100;
            14'h3ff7: o_data_a = 16'b1110110000010000;
            14'h3ff8: o_data_a = 16'b0000000000001101;
            14'h3ff9: o_data_a = 16'b1110001100001000;
            14'h3ffa: o_data_a = 16'b0100010110110011;
            14'h3ffb: o_data_a = 16'b1110110000010000;
            14'h3ffc: o_data_a = 16'b0000000000001110;
            14'h3ffd: o_data_a = 16'b1110001100001000;
            14'h3ffe: o_data_a = 16'b0100000000000010;
            14'h3fff: o_data_a = 16'b1110110000010000;
            14'h4000: o_data_a = 16'b0000000001011111;
            14'h4001: o_data_a = 16'b1110101010000111;
            14'h4002: o_data_a = 16'b0000000000000000;
            14'h4003: o_data_a = 16'b1111110010101000;
            14'h4004: o_data_a = 16'b1111110000010000;
            14'h4005: o_data_a = 16'b0000000000000101;
            14'h4006: o_data_a = 16'b1110001100001000;
            14'h4007: o_data_a = 16'b0000000001101101;
            14'h4008: o_data_a = 16'b1110110000010000;
            14'h4009: o_data_a = 16'b0000000000000000;
            14'h400a: o_data_a = 16'b1111110111101000;
            14'h400b: o_data_a = 16'b1110110010100000;
            14'h400c: o_data_a = 16'b1110001100001000;
            14'h400d: o_data_a = 16'b0000000000000000;
            14'h400e: o_data_a = 16'b1111110111001000;
            14'h400f: o_data_a = 16'b1111110010100000;
            14'h4010: o_data_a = 16'b1110101010001000;
            14'h4011: o_data_a = 16'b0000000000000000;
            14'h4012: o_data_a = 16'b1111110111001000;
            14'h4013: o_data_a = 16'b1111110010100000;
            14'h4014: o_data_a = 16'b1110101010001000;
            14'h4015: o_data_a = 16'b0000000000000000;
            14'h4016: o_data_a = 16'b1111110111001000;
            14'h4017: o_data_a = 16'b1111110010100000;
            14'h4018: o_data_a = 16'b1110101010001000;
            14'h4019: o_data_a = 16'b0000000000011101;
            14'h401a: o_data_a = 16'b1110110000010000;
            14'h401b: o_data_a = 16'b0000000000000000;
            14'h401c: o_data_a = 16'b1111110111101000;
            14'h401d: o_data_a = 16'b1110110010100000;
            14'h401e: o_data_a = 16'b1110001100001000;
            14'h401f: o_data_a = 16'b0000000000111111;
            14'h4020: o_data_a = 16'b1110110000010000;
            14'h4021: o_data_a = 16'b0000000000000000;
            14'h4022: o_data_a = 16'b1111110111101000;
            14'h4023: o_data_a = 16'b1110110010100000;
            14'h4024: o_data_a = 16'b1110001100001000;
            14'h4025: o_data_a = 16'b0000000000101011;
            14'h4026: o_data_a = 16'b1110110000010000;
            14'h4027: o_data_a = 16'b0000000000000000;
            14'h4028: o_data_a = 16'b1111110111101000;
            14'h4029: o_data_a = 16'b1110110010100000;
            14'h402a: o_data_a = 16'b1110001100001000;
            14'h402b: o_data_a = 16'b0000000000101011;
            14'h402c: o_data_a = 16'b1110110000010000;
            14'h402d: o_data_a = 16'b0000000000000000;
            14'h402e: o_data_a = 16'b1111110111101000;
            14'h402f: o_data_a = 16'b1110110010100000;
            14'h4030: o_data_a = 16'b1110001100001000;
            14'h4031: o_data_a = 16'b0000000000101011;
            14'h4032: o_data_a = 16'b1110110000010000;
            14'h4033: o_data_a = 16'b0000000000000000;
            14'h4034: o_data_a = 16'b1111110111101000;
            14'h4035: o_data_a = 16'b1110110010100000;
            14'h4036: o_data_a = 16'b1110001100001000;
            14'h4037: o_data_a = 16'b0000000000101011;
            14'h4038: o_data_a = 16'b1110110000010000;
            14'h4039: o_data_a = 16'b0000000000000000;
            14'h403a: o_data_a = 16'b1111110111101000;
            14'h403b: o_data_a = 16'b1110110010100000;
            14'h403c: o_data_a = 16'b1110001100001000;
            14'h403d: o_data_a = 16'b0000000000000000;
            14'h403e: o_data_a = 16'b1111110111001000;
            14'h403f: o_data_a = 16'b1111110010100000;
            14'h4040: o_data_a = 16'b1110101010001000;
            14'h4041: o_data_a = 16'b0000000000000000;
            14'h4042: o_data_a = 16'b1111110111001000;
            14'h4043: o_data_a = 16'b1111110010100000;
            14'h4044: o_data_a = 16'b1110101010001000;
            14'h4045: o_data_a = 16'b0000000000001100;
            14'h4046: o_data_a = 16'b1110110000010000;
            14'h4047: o_data_a = 16'b0000000000001101;
            14'h4048: o_data_a = 16'b1110001100001000;
            14'h4049: o_data_a = 16'b0100010110110011;
            14'h404a: o_data_a = 16'b1110110000010000;
            14'h404b: o_data_a = 16'b0000000000001110;
            14'h404c: o_data_a = 16'b1110001100001000;
            14'h404d: o_data_a = 16'b0100000001010001;
            14'h404e: o_data_a = 16'b1110110000010000;
            14'h404f: o_data_a = 16'b0000000001011111;
            14'h4050: o_data_a = 16'b1110101010000111;
            14'h4051: o_data_a = 16'b0000000000000000;
            14'h4052: o_data_a = 16'b1111110010101000;
            14'h4053: o_data_a = 16'b1111110000010000;
            14'h4054: o_data_a = 16'b0000000000000101;
            14'h4055: o_data_a = 16'b1110001100001000;
            14'h4056: o_data_a = 16'b0000000001101110;
            14'h4057: o_data_a = 16'b1110110000010000;
            14'h4058: o_data_a = 16'b0000000000000000;
            14'h4059: o_data_a = 16'b1111110111101000;
            14'h405a: o_data_a = 16'b1110110010100000;
            14'h405b: o_data_a = 16'b1110001100001000;
            14'h405c: o_data_a = 16'b0000000000000000;
            14'h405d: o_data_a = 16'b1111110111001000;
            14'h405e: o_data_a = 16'b1111110010100000;
            14'h405f: o_data_a = 16'b1110101010001000;
            14'h4060: o_data_a = 16'b0000000000000000;
            14'h4061: o_data_a = 16'b1111110111001000;
            14'h4062: o_data_a = 16'b1111110010100000;
            14'h4063: o_data_a = 16'b1110101010001000;
            14'h4064: o_data_a = 16'b0000000000000000;
            14'h4065: o_data_a = 16'b1111110111001000;
            14'h4066: o_data_a = 16'b1111110010100000;
            14'h4067: o_data_a = 16'b1110101010001000;
            14'h4068: o_data_a = 16'b0000000000011101;
            14'h4069: o_data_a = 16'b1110110000010000;
            14'h406a: o_data_a = 16'b0000000000000000;
            14'h406b: o_data_a = 16'b1111110111101000;
            14'h406c: o_data_a = 16'b1110110010100000;
            14'h406d: o_data_a = 16'b1110001100001000;
            14'h406e: o_data_a = 16'b0000000000110011;
            14'h406f: o_data_a = 16'b1110110000010000;
            14'h4070: o_data_a = 16'b0000000000000000;
            14'h4071: o_data_a = 16'b1111110111101000;
            14'h4072: o_data_a = 16'b1110110010100000;
            14'h4073: o_data_a = 16'b1110001100001000;
            14'h4074: o_data_a = 16'b0000000000110011;
            14'h4075: o_data_a = 16'b1110110000010000;
            14'h4076: o_data_a = 16'b0000000000000000;
            14'h4077: o_data_a = 16'b1111110111101000;
            14'h4078: o_data_a = 16'b1110110010100000;
            14'h4079: o_data_a = 16'b1110001100001000;
            14'h407a: o_data_a = 16'b0000000000110011;
            14'h407b: o_data_a = 16'b1110110000010000;
            14'h407c: o_data_a = 16'b0000000000000000;
            14'h407d: o_data_a = 16'b1111110111101000;
            14'h407e: o_data_a = 16'b1110110010100000;
            14'h407f: o_data_a = 16'b1110001100001000;
            14'h4080: o_data_a = 16'b0000000000110011;
            14'h4081: o_data_a = 16'b1110110000010000;
            14'h4082: o_data_a = 16'b0000000000000000;
            14'h4083: o_data_a = 16'b1111110111101000;
            14'h4084: o_data_a = 16'b1110110010100000;
            14'h4085: o_data_a = 16'b1110001100001000;
            14'h4086: o_data_a = 16'b0000000000110011;
            14'h4087: o_data_a = 16'b1110110000010000;
            14'h4088: o_data_a = 16'b0000000000000000;
            14'h4089: o_data_a = 16'b1111110111101000;
            14'h408a: o_data_a = 16'b1110110010100000;
            14'h408b: o_data_a = 16'b1110001100001000;
            14'h408c: o_data_a = 16'b0000000000000000;
            14'h408d: o_data_a = 16'b1111110111001000;
            14'h408e: o_data_a = 16'b1111110010100000;
            14'h408f: o_data_a = 16'b1110101010001000;
            14'h4090: o_data_a = 16'b0000000000000000;
            14'h4091: o_data_a = 16'b1111110111001000;
            14'h4092: o_data_a = 16'b1111110010100000;
            14'h4093: o_data_a = 16'b1110101010001000;
            14'h4094: o_data_a = 16'b0000000000001100;
            14'h4095: o_data_a = 16'b1110110000010000;
            14'h4096: o_data_a = 16'b0000000000001101;
            14'h4097: o_data_a = 16'b1110001100001000;
            14'h4098: o_data_a = 16'b0100010110110011;
            14'h4099: o_data_a = 16'b1110110000010000;
            14'h409a: o_data_a = 16'b0000000000001110;
            14'h409b: o_data_a = 16'b1110001100001000;
            14'h409c: o_data_a = 16'b0100000010100000;
            14'h409d: o_data_a = 16'b1110110000010000;
            14'h409e: o_data_a = 16'b0000000001011111;
            14'h409f: o_data_a = 16'b1110101010000111;
            14'h40a0: o_data_a = 16'b0000000000000000;
            14'h40a1: o_data_a = 16'b1111110010101000;
            14'h40a2: o_data_a = 16'b1111110000010000;
            14'h40a3: o_data_a = 16'b0000000000000101;
            14'h40a4: o_data_a = 16'b1110001100001000;
            14'h40a5: o_data_a = 16'b0000000001101111;
            14'h40a6: o_data_a = 16'b1110110000010000;
            14'h40a7: o_data_a = 16'b0000000000000000;
            14'h40a8: o_data_a = 16'b1111110111101000;
            14'h40a9: o_data_a = 16'b1110110010100000;
            14'h40aa: o_data_a = 16'b1110001100001000;
            14'h40ab: o_data_a = 16'b0000000000000000;
            14'h40ac: o_data_a = 16'b1111110111001000;
            14'h40ad: o_data_a = 16'b1111110010100000;
            14'h40ae: o_data_a = 16'b1110101010001000;
            14'h40af: o_data_a = 16'b0000000000000000;
            14'h40b0: o_data_a = 16'b1111110111001000;
            14'h40b1: o_data_a = 16'b1111110010100000;
            14'h40b2: o_data_a = 16'b1110101010001000;
            14'h40b3: o_data_a = 16'b0000000000000000;
            14'h40b4: o_data_a = 16'b1111110111001000;
            14'h40b5: o_data_a = 16'b1111110010100000;
            14'h40b6: o_data_a = 16'b1110101010001000;
            14'h40b7: o_data_a = 16'b0000000000011110;
            14'h40b8: o_data_a = 16'b1110110000010000;
            14'h40b9: o_data_a = 16'b0000000000000000;
            14'h40ba: o_data_a = 16'b1111110111101000;
            14'h40bb: o_data_a = 16'b1110110010100000;
            14'h40bc: o_data_a = 16'b1110001100001000;
            14'h40bd: o_data_a = 16'b0000000000110011;
            14'h40be: o_data_a = 16'b1110110000010000;
            14'h40bf: o_data_a = 16'b0000000000000000;
            14'h40c0: o_data_a = 16'b1111110111101000;
            14'h40c1: o_data_a = 16'b1110110010100000;
            14'h40c2: o_data_a = 16'b1110001100001000;
            14'h40c3: o_data_a = 16'b0000000000110011;
            14'h40c4: o_data_a = 16'b1110110000010000;
            14'h40c5: o_data_a = 16'b0000000000000000;
            14'h40c6: o_data_a = 16'b1111110111101000;
            14'h40c7: o_data_a = 16'b1110110010100000;
            14'h40c8: o_data_a = 16'b1110001100001000;
            14'h40c9: o_data_a = 16'b0000000000110011;
            14'h40ca: o_data_a = 16'b1110110000010000;
            14'h40cb: o_data_a = 16'b0000000000000000;
            14'h40cc: o_data_a = 16'b1111110111101000;
            14'h40cd: o_data_a = 16'b1110110010100000;
            14'h40ce: o_data_a = 16'b1110001100001000;
            14'h40cf: o_data_a = 16'b0000000000110011;
            14'h40d0: o_data_a = 16'b1110110000010000;
            14'h40d1: o_data_a = 16'b0000000000000000;
            14'h40d2: o_data_a = 16'b1111110111101000;
            14'h40d3: o_data_a = 16'b1110110010100000;
            14'h40d4: o_data_a = 16'b1110001100001000;
            14'h40d5: o_data_a = 16'b0000000000011110;
            14'h40d6: o_data_a = 16'b1110110000010000;
            14'h40d7: o_data_a = 16'b0000000000000000;
            14'h40d8: o_data_a = 16'b1111110111101000;
            14'h40d9: o_data_a = 16'b1110110010100000;
            14'h40da: o_data_a = 16'b1110001100001000;
            14'h40db: o_data_a = 16'b0000000000000000;
            14'h40dc: o_data_a = 16'b1111110111001000;
            14'h40dd: o_data_a = 16'b1111110010100000;
            14'h40de: o_data_a = 16'b1110101010001000;
            14'h40df: o_data_a = 16'b0000000000000000;
            14'h40e0: o_data_a = 16'b1111110111001000;
            14'h40e1: o_data_a = 16'b1111110010100000;
            14'h40e2: o_data_a = 16'b1110101010001000;
            14'h40e3: o_data_a = 16'b0000000000001100;
            14'h40e4: o_data_a = 16'b1110110000010000;
            14'h40e5: o_data_a = 16'b0000000000001101;
            14'h40e6: o_data_a = 16'b1110001100001000;
            14'h40e7: o_data_a = 16'b0100010110110011;
            14'h40e8: o_data_a = 16'b1110110000010000;
            14'h40e9: o_data_a = 16'b0000000000001110;
            14'h40ea: o_data_a = 16'b1110001100001000;
            14'h40eb: o_data_a = 16'b0100000011101111;
            14'h40ec: o_data_a = 16'b1110110000010000;
            14'h40ed: o_data_a = 16'b0000000001011111;
            14'h40ee: o_data_a = 16'b1110101010000111;
            14'h40ef: o_data_a = 16'b0000000000000000;
            14'h40f0: o_data_a = 16'b1111110010101000;
            14'h40f1: o_data_a = 16'b1111110000010000;
            14'h40f2: o_data_a = 16'b0000000000000101;
            14'h40f3: o_data_a = 16'b1110001100001000;
            14'h40f4: o_data_a = 16'b0000000001110000;
            14'h40f5: o_data_a = 16'b1110110000010000;
            14'h40f6: o_data_a = 16'b0000000000000000;
            14'h40f7: o_data_a = 16'b1111110111101000;
            14'h40f8: o_data_a = 16'b1110110010100000;
            14'h40f9: o_data_a = 16'b1110001100001000;
            14'h40fa: o_data_a = 16'b0000000000000000;
            14'h40fb: o_data_a = 16'b1111110111001000;
            14'h40fc: o_data_a = 16'b1111110010100000;
            14'h40fd: o_data_a = 16'b1110101010001000;
            14'h40fe: o_data_a = 16'b0000000000000000;
            14'h40ff: o_data_a = 16'b1111110111001000;
            14'h4100: o_data_a = 16'b1111110010100000;
            14'h4101: o_data_a = 16'b1110101010001000;
            14'h4102: o_data_a = 16'b0000000000000000;
            14'h4103: o_data_a = 16'b1111110111001000;
            14'h4104: o_data_a = 16'b1111110010100000;
            14'h4105: o_data_a = 16'b1110101010001000;
            14'h4106: o_data_a = 16'b0000000000011110;
            14'h4107: o_data_a = 16'b1110110000010000;
            14'h4108: o_data_a = 16'b0000000000000000;
            14'h4109: o_data_a = 16'b1111110111101000;
            14'h410a: o_data_a = 16'b1110110010100000;
            14'h410b: o_data_a = 16'b1110001100001000;
            14'h410c: o_data_a = 16'b0000000000110011;
            14'h410d: o_data_a = 16'b1110110000010000;
            14'h410e: o_data_a = 16'b0000000000000000;
            14'h410f: o_data_a = 16'b1111110111101000;
            14'h4110: o_data_a = 16'b1110110010100000;
            14'h4111: o_data_a = 16'b1110001100001000;
            14'h4112: o_data_a = 16'b0000000000110011;
            14'h4113: o_data_a = 16'b1110110000010000;
            14'h4114: o_data_a = 16'b0000000000000000;
            14'h4115: o_data_a = 16'b1111110111101000;
            14'h4116: o_data_a = 16'b1110110010100000;
            14'h4117: o_data_a = 16'b1110001100001000;
            14'h4118: o_data_a = 16'b0000000000110011;
            14'h4119: o_data_a = 16'b1110110000010000;
            14'h411a: o_data_a = 16'b0000000000000000;
            14'h411b: o_data_a = 16'b1111110111101000;
            14'h411c: o_data_a = 16'b1110110010100000;
            14'h411d: o_data_a = 16'b1110001100001000;
            14'h411e: o_data_a = 16'b0000000000011111;
            14'h411f: o_data_a = 16'b1110110000010000;
            14'h4120: o_data_a = 16'b0000000000000000;
            14'h4121: o_data_a = 16'b1111110111101000;
            14'h4122: o_data_a = 16'b1110110010100000;
            14'h4123: o_data_a = 16'b1110001100001000;
            14'h4124: o_data_a = 16'b0000000000000011;
            14'h4125: o_data_a = 16'b1110110000010000;
            14'h4126: o_data_a = 16'b0000000000000000;
            14'h4127: o_data_a = 16'b1111110111101000;
            14'h4128: o_data_a = 16'b1110110010100000;
            14'h4129: o_data_a = 16'b1110001100001000;
            14'h412a: o_data_a = 16'b0000000000000011;
            14'h412b: o_data_a = 16'b1110110000010000;
            14'h412c: o_data_a = 16'b0000000000000000;
            14'h412d: o_data_a = 16'b1111110111101000;
            14'h412e: o_data_a = 16'b1110110010100000;
            14'h412f: o_data_a = 16'b1110001100001000;
            14'h4130: o_data_a = 16'b0000000000000000;
            14'h4131: o_data_a = 16'b1111110111001000;
            14'h4132: o_data_a = 16'b1111110010100000;
            14'h4133: o_data_a = 16'b1110101010001000;
            14'h4134: o_data_a = 16'b0000000000001100;
            14'h4135: o_data_a = 16'b1110110000010000;
            14'h4136: o_data_a = 16'b0000000000001101;
            14'h4137: o_data_a = 16'b1110001100001000;
            14'h4138: o_data_a = 16'b0100010110110011;
            14'h4139: o_data_a = 16'b1110110000010000;
            14'h413a: o_data_a = 16'b0000000000001110;
            14'h413b: o_data_a = 16'b1110001100001000;
            14'h413c: o_data_a = 16'b0100000101000000;
            14'h413d: o_data_a = 16'b1110110000010000;
            14'h413e: o_data_a = 16'b0000000001011111;
            14'h413f: o_data_a = 16'b1110101010000111;
            14'h4140: o_data_a = 16'b0000000000000000;
            14'h4141: o_data_a = 16'b1111110010101000;
            14'h4142: o_data_a = 16'b1111110000010000;
            14'h4143: o_data_a = 16'b0000000000000101;
            14'h4144: o_data_a = 16'b1110001100001000;
            14'h4145: o_data_a = 16'b0000000001110001;
            14'h4146: o_data_a = 16'b1110110000010000;
            14'h4147: o_data_a = 16'b0000000000000000;
            14'h4148: o_data_a = 16'b1111110111101000;
            14'h4149: o_data_a = 16'b1110110010100000;
            14'h414a: o_data_a = 16'b1110001100001000;
            14'h414b: o_data_a = 16'b0000000000000000;
            14'h414c: o_data_a = 16'b1111110111001000;
            14'h414d: o_data_a = 16'b1111110010100000;
            14'h414e: o_data_a = 16'b1110101010001000;
            14'h414f: o_data_a = 16'b0000000000000000;
            14'h4150: o_data_a = 16'b1111110111001000;
            14'h4151: o_data_a = 16'b1111110010100000;
            14'h4152: o_data_a = 16'b1110101010001000;
            14'h4153: o_data_a = 16'b0000000000000000;
            14'h4154: o_data_a = 16'b1111110111001000;
            14'h4155: o_data_a = 16'b1111110010100000;
            14'h4156: o_data_a = 16'b1110101010001000;
            14'h4157: o_data_a = 16'b0000000000011110;
            14'h4158: o_data_a = 16'b1110110000010000;
            14'h4159: o_data_a = 16'b0000000000000000;
            14'h415a: o_data_a = 16'b1111110111101000;
            14'h415b: o_data_a = 16'b1110110010100000;
            14'h415c: o_data_a = 16'b1110001100001000;
            14'h415d: o_data_a = 16'b0000000000110011;
            14'h415e: o_data_a = 16'b1110110000010000;
            14'h415f: o_data_a = 16'b0000000000000000;
            14'h4160: o_data_a = 16'b1111110111101000;
            14'h4161: o_data_a = 16'b1110110010100000;
            14'h4162: o_data_a = 16'b1110001100001000;
            14'h4163: o_data_a = 16'b0000000000110011;
            14'h4164: o_data_a = 16'b1110110000010000;
            14'h4165: o_data_a = 16'b0000000000000000;
            14'h4166: o_data_a = 16'b1111110111101000;
            14'h4167: o_data_a = 16'b1110110010100000;
            14'h4168: o_data_a = 16'b1110001100001000;
            14'h4169: o_data_a = 16'b0000000000110011;
            14'h416a: o_data_a = 16'b1110110000010000;
            14'h416b: o_data_a = 16'b0000000000000000;
            14'h416c: o_data_a = 16'b1111110111101000;
            14'h416d: o_data_a = 16'b1110110010100000;
            14'h416e: o_data_a = 16'b1110001100001000;
            14'h416f: o_data_a = 16'b0000000000111110;
            14'h4170: o_data_a = 16'b1110110000010000;
            14'h4171: o_data_a = 16'b0000000000000000;
            14'h4172: o_data_a = 16'b1111110111101000;
            14'h4173: o_data_a = 16'b1110110010100000;
            14'h4174: o_data_a = 16'b1110001100001000;
            14'h4175: o_data_a = 16'b0000000000110000;
            14'h4176: o_data_a = 16'b1110110000010000;
            14'h4177: o_data_a = 16'b0000000000000000;
            14'h4178: o_data_a = 16'b1111110111101000;
            14'h4179: o_data_a = 16'b1110110010100000;
            14'h417a: o_data_a = 16'b1110001100001000;
            14'h417b: o_data_a = 16'b0000000000110000;
            14'h417c: o_data_a = 16'b1110110000010000;
            14'h417d: o_data_a = 16'b0000000000000000;
            14'h417e: o_data_a = 16'b1111110111101000;
            14'h417f: o_data_a = 16'b1110110010100000;
            14'h4180: o_data_a = 16'b1110001100001000;
            14'h4181: o_data_a = 16'b0000000000000000;
            14'h4182: o_data_a = 16'b1111110111001000;
            14'h4183: o_data_a = 16'b1111110010100000;
            14'h4184: o_data_a = 16'b1110101010001000;
            14'h4185: o_data_a = 16'b0000000000001100;
            14'h4186: o_data_a = 16'b1110110000010000;
            14'h4187: o_data_a = 16'b0000000000001101;
            14'h4188: o_data_a = 16'b1110001100001000;
            14'h4189: o_data_a = 16'b0100010110110011;
            14'h418a: o_data_a = 16'b1110110000010000;
            14'h418b: o_data_a = 16'b0000000000001110;
            14'h418c: o_data_a = 16'b1110001100001000;
            14'h418d: o_data_a = 16'b0100000110010001;
            14'h418e: o_data_a = 16'b1110110000010000;
            14'h418f: o_data_a = 16'b0000000001011111;
            14'h4190: o_data_a = 16'b1110101010000111;
            14'h4191: o_data_a = 16'b0000000000000000;
            14'h4192: o_data_a = 16'b1111110010101000;
            14'h4193: o_data_a = 16'b1111110000010000;
            14'h4194: o_data_a = 16'b0000000000000101;
            14'h4195: o_data_a = 16'b1110001100001000;
            14'h4196: o_data_a = 16'b0000000001110010;
            14'h4197: o_data_a = 16'b1110110000010000;
            14'h4198: o_data_a = 16'b0000000000000000;
            14'h4199: o_data_a = 16'b1111110111101000;
            14'h419a: o_data_a = 16'b1110110010100000;
            14'h419b: o_data_a = 16'b1110001100001000;
            14'h419c: o_data_a = 16'b0000000000000000;
            14'h419d: o_data_a = 16'b1111110111001000;
            14'h419e: o_data_a = 16'b1111110010100000;
            14'h419f: o_data_a = 16'b1110101010001000;
            14'h41a0: o_data_a = 16'b0000000000000000;
            14'h41a1: o_data_a = 16'b1111110111001000;
            14'h41a2: o_data_a = 16'b1111110010100000;
            14'h41a3: o_data_a = 16'b1110101010001000;
            14'h41a4: o_data_a = 16'b0000000000000000;
            14'h41a5: o_data_a = 16'b1111110111001000;
            14'h41a6: o_data_a = 16'b1111110010100000;
            14'h41a7: o_data_a = 16'b1110101010001000;
            14'h41a8: o_data_a = 16'b0000000000011101;
            14'h41a9: o_data_a = 16'b1110110000010000;
            14'h41aa: o_data_a = 16'b0000000000000000;
            14'h41ab: o_data_a = 16'b1111110111101000;
            14'h41ac: o_data_a = 16'b1110110010100000;
            14'h41ad: o_data_a = 16'b1110001100001000;
            14'h41ae: o_data_a = 16'b0000000000110111;
            14'h41af: o_data_a = 16'b1110110000010000;
            14'h41b0: o_data_a = 16'b0000000000000000;
            14'h41b1: o_data_a = 16'b1111110111101000;
            14'h41b2: o_data_a = 16'b1110110010100000;
            14'h41b3: o_data_a = 16'b1110001100001000;
            14'h41b4: o_data_a = 16'b0000000000110011;
            14'h41b5: o_data_a = 16'b1110110000010000;
            14'h41b6: o_data_a = 16'b0000000000000000;
            14'h41b7: o_data_a = 16'b1111110111101000;
            14'h41b8: o_data_a = 16'b1110110010100000;
            14'h41b9: o_data_a = 16'b1110001100001000;
            14'h41ba: o_data_a = 16'b0000000000000011;
            14'h41bb: o_data_a = 16'b1110110000010000;
            14'h41bc: o_data_a = 16'b0000000000000000;
            14'h41bd: o_data_a = 16'b1111110111101000;
            14'h41be: o_data_a = 16'b1110110010100000;
            14'h41bf: o_data_a = 16'b1110001100001000;
            14'h41c0: o_data_a = 16'b0000000000000011;
            14'h41c1: o_data_a = 16'b1110110000010000;
            14'h41c2: o_data_a = 16'b0000000000000000;
            14'h41c3: o_data_a = 16'b1111110111101000;
            14'h41c4: o_data_a = 16'b1110110010100000;
            14'h41c5: o_data_a = 16'b1110001100001000;
            14'h41c6: o_data_a = 16'b0000000000000111;
            14'h41c7: o_data_a = 16'b1110110000010000;
            14'h41c8: o_data_a = 16'b0000000000000000;
            14'h41c9: o_data_a = 16'b1111110111101000;
            14'h41ca: o_data_a = 16'b1110110010100000;
            14'h41cb: o_data_a = 16'b1110001100001000;
            14'h41cc: o_data_a = 16'b0000000000000000;
            14'h41cd: o_data_a = 16'b1111110111001000;
            14'h41ce: o_data_a = 16'b1111110010100000;
            14'h41cf: o_data_a = 16'b1110101010001000;
            14'h41d0: o_data_a = 16'b0000000000000000;
            14'h41d1: o_data_a = 16'b1111110111001000;
            14'h41d2: o_data_a = 16'b1111110010100000;
            14'h41d3: o_data_a = 16'b1110101010001000;
            14'h41d4: o_data_a = 16'b0000000000001100;
            14'h41d5: o_data_a = 16'b1110110000010000;
            14'h41d6: o_data_a = 16'b0000000000001101;
            14'h41d7: o_data_a = 16'b1110001100001000;
            14'h41d8: o_data_a = 16'b0100010110110011;
            14'h41d9: o_data_a = 16'b1110110000010000;
            14'h41da: o_data_a = 16'b0000000000001110;
            14'h41db: o_data_a = 16'b1110001100001000;
            14'h41dc: o_data_a = 16'b0100000111100000;
            14'h41dd: o_data_a = 16'b1110110000010000;
            14'h41de: o_data_a = 16'b0000000001011111;
            14'h41df: o_data_a = 16'b1110101010000111;
            14'h41e0: o_data_a = 16'b0000000000000000;
            14'h41e1: o_data_a = 16'b1111110010101000;
            14'h41e2: o_data_a = 16'b1111110000010000;
            14'h41e3: o_data_a = 16'b0000000000000101;
            14'h41e4: o_data_a = 16'b1110001100001000;
            14'h41e5: o_data_a = 16'b0000000001110011;
            14'h41e6: o_data_a = 16'b1110110000010000;
            14'h41e7: o_data_a = 16'b0000000000000000;
            14'h41e8: o_data_a = 16'b1111110111101000;
            14'h41e9: o_data_a = 16'b1110110010100000;
            14'h41ea: o_data_a = 16'b1110001100001000;
            14'h41eb: o_data_a = 16'b0000000000000000;
            14'h41ec: o_data_a = 16'b1111110111001000;
            14'h41ed: o_data_a = 16'b1111110010100000;
            14'h41ee: o_data_a = 16'b1110101010001000;
            14'h41ef: o_data_a = 16'b0000000000000000;
            14'h41f0: o_data_a = 16'b1111110111001000;
            14'h41f1: o_data_a = 16'b1111110010100000;
            14'h41f2: o_data_a = 16'b1110101010001000;
            14'h41f3: o_data_a = 16'b0000000000000000;
            14'h41f4: o_data_a = 16'b1111110111001000;
            14'h41f5: o_data_a = 16'b1111110010100000;
            14'h41f6: o_data_a = 16'b1110101010001000;
            14'h41f7: o_data_a = 16'b0000000000011110;
            14'h41f8: o_data_a = 16'b1110110000010000;
            14'h41f9: o_data_a = 16'b0000000000000000;
            14'h41fa: o_data_a = 16'b1111110111101000;
            14'h41fb: o_data_a = 16'b1110110010100000;
            14'h41fc: o_data_a = 16'b1110001100001000;
            14'h41fd: o_data_a = 16'b0000000000110011;
            14'h41fe: o_data_a = 16'b1110110000010000;
            14'h41ff: o_data_a = 16'b0000000000000000;
            14'h4200: o_data_a = 16'b1111110111101000;
            14'h4201: o_data_a = 16'b1110110010100000;
            14'h4202: o_data_a = 16'b1110001100001000;
            14'h4203: o_data_a = 16'b0000000000000110;
            14'h4204: o_data_a = 16'b1110110000010000;
            14'h4205: o_data_a = 16'b0000000000000000;
            14'h4206: o_data_a = 16'b1111110111101000;
            14'h4207: o_data_a = 16'b1110110010100000;
            14'h4208: o_data_a = 16'b1110001100001000;
            14'h4209: o_data_a = 16'b0000000000011000;
            14'h420a: o_data_a = 16'b1110110000010000;
            14'h420b: o_data_a = 16'b0000000000000000;
            14'h420c: o_data_a = 16'b1111110111101000;
            14'h420d: o_data_a = 16'b1110110010100000;
            14'h420e: o_data_a = 16'b1110001100001000;
            14'h420f: o_data_a = 16'b0000000000110011;
            14'h4210: o_data_a = 16'b1110110000010000;
            14'h4211: o_data_a = 16'b0000000000000000;
            14'h4212: o_data_a = 16'b1111110111101000;
            14'h4213: o_data_a = 16'b1110110010100000;
            14'h4214: o_data_a = 16'b1110001100001000;
            14'h4215: o_data_a = 16'b0000000000011110;
            14'h4216: o_data_a = 16'b1110110000010000;
            14'h4217: o_data_a = 16'b0000000000000000;
            14'h4218: o_data_a = 16'b1111110111101000;
            14'h4219: o_data_a = 16'b1110110010100000;
            14'h421a: o_data_a = 16'b1110001100001000;
            14'h421b: o_data_a = 16'b0000000000000000;
            14'h421c: o_data_a = 16'b1111110111001000;
            14'h421d: o_data_a = 16'b1111110010100000;
            14'h421e: o_data_a = 16'b1110101010001000;
            14'h421f: o_data_a = 16'b0000000000000000;
            14'h4220: o_data_a = 16'b1111110111001000;
            14'h4221: o_data_a = 16'b1111110010100000;
            14'h4222: o_data_a = 16'b1110101010001000;
            14'h4223: o_data_a = 16'b0000000000001100;
            14'h4224: o_data_a = 16'b1110110000010000;
            14'h4225: o_data_a = 16'b0000000000001101;
            14'h4226: o_data_a = 16'b1110001100001000;
            14'h4227: o_data_a = 16'b0100010110110011;
            14'h4228: o_data_a = 16'b1110110000010000;
            14'h4229: o_data_a = 16'b0000000000001110;
            14'h422a: o_data_a = 16'b1110001100001000;
            14'h422b: o_data_a = 16'b0100001000101111;
            14'h422c: o_data_a = 16'b1110110000010000;
            14'h422d: o_data_a = 16'b0000000001011111;
            14'h422e: o_data_a = 16'b1110101010000111;
            14'h422f: o_data_a = 16'b0000000000000000;
            14'h4230: o_data_a = 16'b1111110010101000;
            14'h4231: o_data_a = 16'b1111110000010000;
            14'h4232: o_data_a = 16'b0000000000000101;
            14'h4233: o_data_a = 16'b1110001100001000;
            14'h4234: o_data_a = 16'b0000000001110100;
            14'h4235: o_data_a = 16'b1110110000010000;
            14'h4236: o_data_a = 16'b0000000000000000;
            14'h4237: o_data_a = 16'b1111110111101000;
            14'h4238: o_data_a = 16'b1110110010100000;
            14'h4239: o_data_a = 16'b1110001100001000;
            14'h423a: o_data_a = 16'b0000000000000100;
            14'h423b: o_data_a = 16'b1110110000010000;
            14'h423c: o_data_a = 16'b0000000000000000;
            14'h423d: o_data_a = 16'b1111110111101000;
            14'h423e: o_data_a = 16'b1110110010100000;
            14'h423f: o_data_a = 16'b1110001100001000;
            14'h4240: o_data_a = 16'b0000000000000110;
            14'h4241: o_data_a = 16'b1110110000010000;
            14'h4242: o_data_a = 16'b0000000000000000;
            14'h4243: o_data_a = 16'b1111110111101000;
            14'h4244: o_data_a = 16'b1110110010100000;
            14'h4245: o_data_a = 16'b1110001100001000;
            14'h4246: o_data_a = 16'b0000000000000110;
            14'h4247: o_data_a = 16'b1110110000010000;
            14'h4248: o_data_a = 16'b0000000000000000;
            14'h4249: o_data_a = 16'b1111110111101000;
            14'h424a: o_data_a = 16'b1110110010100000;
            14'h424b: o_data_a = 16'b1110001100001000;
            14'h424c: o_data_a = 16'b0000000000001111;
            14'h424d: o_data_a = 16'b1110110000010000;
            14'h424e: o_data_a = 16'b0000000000000000;
            14'h424f: o_data_a = 16'b1111110111101000;
            14'h4250: o_data_a = 16'b1110110010100000;
            14'h4251: o_data_a = 16'b1110001100001000;
            14'h4252: o_data_a = 16'b0000000000000110;
            14'h4253: o_data_a = 16'b1110110000010000;
            14'h4254: o_data_a = 16'b0000000000000000;
            14'h4255: o_data_a = 16'b1111110111101000;
            14'h4256: o_data_a = 16'b1110110010100000;
            14'h4257: o_data_a = 16'b1110001100001000;
            14'h4258: o_data_a = 16'b0000000000000110;
            14'h4259: o_data_a = 16'b1110110000010000;
            14'h425a: o_data_a = 16'b0000000000000000;
            14'h425b: o_data_a = 16'b1111110111101000;
            14'h425c: o_data_a = 16'b1110110010100000;
            14'h425d: o_data_a = 16'b1110001100001000;
            14'h425e: o_data_a = 16'b0000000000000110;
            14'h425f: o_data_a = 16'b1110110000010000;
            14'h4260: o_data_a = 16'b0000000000000000;
            14'h4261: o_data_a = 16'b1111110111101000;
            14'h4262: o_data_a = 16'b1110110010100000;
            14'h4263: o_data_a = 16'b1110001100001000;
            14'h4264: o_data_a = 16'b0000000000110110;
            14'h4265: o_data_a = 16'b1110110000010000;
            14'h4266: o_data_a = 16'b0000000000000000;
            14'h4267: o_data_a = 16'b1111110111101000;
            14'h4268: o_data_a = 16'b1110110010100000;
            14'h4269: o_data_a = 16'b1110001100001000;
            14'h426a: o_data_a = 16'b0000000000011100;
            14'h426b: o_data_a = 16'b1110110000010000;
            14'h426c: o_data_a = 16'b0000000000000000;
            14'h426d: o_data_a = 16'b1111110111101000;
            14'h426e: o_data_a = 16'b1110110010100000;
            14'h426f: o_data_a = 16'b1110001100001000;
            14'h4270: o_data_a = 16'b0000000000000000;
            14'h4271: o_data_a = 16'b1111110111001000;
            14'h4272: o_data_a = 16'b1111110010100000;
            14'h4273: o_data_a = 16'b1110101010001000;
            14'h4274: o_data_a = 16'b0000000000000000;
            14'h4275: o_data_a = 16'b1111110111001000;
            14'h4276: o_data_a = 16'b1111110010100000;
            14'h4277: o_data_a = 16'b1110101010001000;
            14'h4278: o_data_a = 16'b0000000000001100;
            14'h4279: o_data_a = 16'b1110110000010000;
            14'h427a: o_data_a = 16'b0000000000001101;
            14'h427b: o_data_a = 16'b1110001100001000;
            14'h427c: o_data_a = 16'b0100010110110011;
            14'h427d: o_data_a = 16'b1110110000010000;
            14'h427e: o_data_a = 16'b0000000000001110;
            14'h427f: o_data_a = 16'b1110001100001000;
            14'h4280: o_data_a = 16'b0100001010000100;
            14'h4281: o_data_a = 16'b1110110000010000;
            14'h4282: o_data_a = 16'b0000000001011111;
            14'h4283: o_data_a = 16'b1110101010000111;
            14'h4284: o_data_a = 16'b0000000000000000;
            14'h4285: o_data_a = 16'b1111110010101000;
            14'h4286: o_data_a = 16'b1111110000010000;
            14'h4287: o_data_a = 16'b0000000000000101;
            14'h4288: o_data_a = 16'b1110001100001000;
            14'h4289: o_data_a = 16'b0000000001110101;
            14'h428a: o_data_a = 16'b1110110000010000;
            14'h428b: o_data_a = 16'b0000000000000000;
            14'h428c: o_data_a = 16'b1111110111101000;
            14'h428d: o_data_a = 16'b1110110010100000;
            14'h428e: o_data_a = 16'b1110001100001000;
            14'h428f: o_data_a = 16'b0000000000000000;
            14'h4290: o_data_a = 16'b1111110111001000;
            14'h4291: o_data_a = 16'b1111110010100000;
            14'h4292: o_data_a = 16'b1110101010001000;
            14'h4293: o_data_a = 16'b0000000000000000;
            14'h4294: o_data_a = 16'b1111110111001000;
            14'h4295: o_data_a = 16'b1111110010100000;
            14'h4296: o_data_a = 16'b1110101010001000;
            14'h4297: o_data_a = 16'b0000000000000000;
            14'h4298: o_data_a = 16'b1111110111001000;
            14'h4299: o_data_a = 16'b1111110010100000;
            14'h429a: o_data_a = 16'b1110101010001000;
            14'h429b: o_data_a = 16'b0000000000011011;
            14'h429c: o_data_a = 16'b1110110000010000;
            14'h429d: o_data_a = 16'b0000000000000000;
            14'h429e: o_data_a = 16'b1111110111101000;
            14'h429f: o_data_a = 16'b1110110010100000;
            14'h42a0: o_data_a = 16'b1110001100001000;
            14'h42a1: o_data_a = 16'b0000000000011011;
            14'h42a2: o_data_a = 16'b1110110000010000;
            14'h42a3: o_data_a = 16'b0000000000000000;
            14'h42a4: o_data_a = 16'b1111110111101000;
            14'h42a5: o_data_a = 16'b1110110010100000;
            14'h42a6: o_data_a = 16'b1110001100001000;
            14'h42a7: o_data_a = 16'b0000000000011011;
            14'h42a8: o_data_a = 16'b1110110000010000;
            14'h42a9: o_data_a = 16'b0000000000000000;
            14'h42aa: o_data_a = 16'b1111110111101000;
            14'h42ab: o_data_a = 16'b1110110010100000;
            14'h42ac: o_data_a = 16'b1110001100001000;
            14'h42ad: o_data_a = 16'b0000000000011011;
            14'h42ae: o_data_a = 16'b1110110000010000;
            14'h42af: o_data_a = 16'b0000000000000000;
            14'h42b0: o_data_a = 16'b1111110111101000;
            14'h42b1: o_data_a = 16'b1110110010100000;
            14'h42b2: o_data_a = 16'b1110001100001000;
            14'h42b3: o_data_a = 16'b0000000000011011;
            14'h42b4: o_data_a = 16'b1110110000010000;
            14'h42b5: o_data_a = 16'b0000000000000000;
            14'h42b6: o_data_a = 16'b1111110111101000;
            14'h42b7: o_data_a = 16'b1110110010100000;
            14'h42b8: o_data_a = 16'b1110001100001000;
            14'h42b9: o_data_a = 16'b0000000000110110;
            14'h42ba: o_data_a = 16'b1110110000010000;
            14'h42bb: o_data_a = 16'b0000000000000000;
            14'h42bc: o_data_a = 16'b1111110111101000;
            14'h42bd: o_data_a = 16'b1110110010100000;
            14'h42be: o_data_a = 16'b1110001100001000;
            14'h42bf: o_data_a = 16'b0000000000000000;
            14'h42c0: o_data_a = 16'b1111110111001000;
            14'h42c1: o_data_a = 16'b1111110010100000;
            14'h42c2: o_data_a = 16'b1110101010001000;
            14'h42c3: o_data_a = 16'b0000000000000000;
            14'h42c4: o_data_a = 16'b1111110111001000;
            14'h42c5: o_data_a = 16'b1111110010100000;
            14'h42c6: o_data_a = 16'b1110101010001000;
            14'h42c7: o_data_a = 16'b0000000000001100;
            14'h42c8: o_data_a = 16'b1110110000010000;
            14'h42c9: o_data_a = 16'b0000000000001101;
            14'h42ca: o_data_a = 16'b1110001100001000;
            14'h42cb: o_data_a = 16'b0100010110110011;
            14'h42cc: o_data_a = 16'b1110110000010000;
            14'h42cd: o_data_a = 16'b0000000000001110;
            14'h42ce: o_data_a = 16'b1110001100001000;
            14'h42cf: o_data_a = 16'b0100001011010011;
            14'h42d0: o_data_a = 16'b1110110000010000;
            14'h42d1: o_data_a = 16'b0000000001011111;
            14'h42d2: o_data_a = 16'b1110101010000111;
            14'h42d3: o_data_a = 16'b0000000000000000;
            14'h42d4: o_data_a = 16'b1111110010101000;
            14'h42d5: o_data_a = 16'b1111110000010000;
            14'h42d6: o_data_a = 16'b0000000000000101;
            14'h42d7: o_data_a = 16'b1110001100001000;
            14'h42d8: o_data_a = 16'b0000000001110110;
            14'h42d9: o_data_a = 16'b1110110000010000;
            14'h42da: o_data_a = 16'b0000000000000000;
            14'h42db: o_data_a = 16'b1111110111101000;
            14'h42dc: o_data_a = 16'b1110110010100000;
            14'h42dd: o_data_a = 16'b1110001100001000;
            14'h42de: o_data_a = 16'b0000000000000000;
            14'h42df: o_data_a = 16'b1111110111001000;
            14'h42e0: o_data_a = 16'b1111110010100000;
            14'h42e1: o_data_a = 16'b1110101010001000;
            14'h42e2: o_data_a = 16'b0000000000000000;
            14'h42e3: o_data_a = 16'b1111110111001000;
            14'h42e4: o_data_a = 16'b1111110010100000;
            14'h42e5: o_data_a = 16'b1110101010001000;
            14'h42e6: o_data_a = 16'b0000000000000000;
            14'h42e7: o_data_a = 16'b1111110111001000;
            14'h42e8: o_data_a = 16'b1111110010100000;
            14'h42e9: o_data_a = 16'b1110101010001000;
            14'h42ea: o_data_a = 16'b0000000000110011;
            14'h42eb: o_data_a = 16'b1110110000010000;
            14'h42ec: o_data_a = 16'b0000000000000000;
            14'h42ed: o_data_a = 16'b1111110111101000;
            14'h42ee: o_data_a = 16'b1110110010100000;
            14'h42ef: o_data_a = 16'b1110001100001000;
            14'h42f0: o_data_a = 16'b0000000000110011;
            14'h42f1: o_data_a = 16'b1110110000010000;
            14'h42f2: o_data_a = 16'b0000000000000000;
            14'h42f3: o_data_a = 16'b1111110111101000;
            14'h42f4: o_data_a = 16'b1110110010100000;
            14'h42f5: o_data_a = 16'b1110001100001000;
            14'h42f6: o_data_a = 16'b0000000000110011;
            14'h42f7: o_data_a = 16'b1110110000010000;
            14'h42f8: o_data_a = 16'b0000000000000000;
            14'h42f9: o_data_a = 16'b1111110111101000;
            14'h42fa: o_data_a = 16'b1110110010100000;
            14'h42fb: o_data_a = 16'b1110001100001000;
            14'h42fc: o_data_a = 16'b0000000000110011;
            14'h42fd: o_data_a = 16'b1110110000010000;
            14'h42fe: o_data_a = 16'b0000000000000000;
            14'h42ff: o_data_a = 16'b1111110111101000;
            14'h4300: o_data_a = 16'b1110110010100000;
            14'h4301: o_data_a = 16'b1110001100001000;
            14'h4302: o_data_a = 16'b0000000000011110;
            14'h4303: o_data_a = 16'b1110110000010000;
            14'h4304: o_data_a = 16'b0000000000000000;
            14'h4305: o_data_a = 16'b1111110111101000;
            14'h4306: o_data_a = 16'b1110110010100000;
            14'h4307: o_data_a = 16'b1110001100001000;
            14'h4308: o_data_a = 16'b0000000000001100;
            14'h4309: o_data_a = 16'b1110110000010000;
            14'h430a: o_data_a = 16'b0000000000000000;
            14'h430b: o_data_a = 16'b1111110111101000;
            14'h430c: o_data_a = 16'b1110110010100000;
            14'h430d: o_data_a = 16'b1110001100001000;
            14'h430e: o_data_a = 16'b0000000000000000;
            14'h430f: o_data_a = 16'b1111110111001000;
            14'h4310: o_data_a = 16'b1111110010100000;
            14'h4311: o_data_a = 16'b1110101010001000;
            14'h4312: o_data_a = 16'b0000000000000000;
            14'h4313: o_data_a = 16'b1111110111001000;
            14'h4314: o_data_a = 16'b1111110010100000;
            14'h4315: o_data_a = 16'b1110101010001000;
            14'h4316: o_data_a = 16'b0000000000001100;
            14'h4317: o_data_a = 16'b1110110000010000;
            14'h4318: o_data_a = 16'b0000000000001101;
            14'h4319: o_data_a = 16'b1110001100001000;
            14'h431a: o_data_a = 16'b0100010110110011;
            14'h431b: o_data_a = 16'b1110110000010000;
            14'h431c: o_data_a = 16'b0000000000001110;
            14'h431d: o_data_a = 16'b1110001100001000;
            14'h431e: o_data_a = 16'b0100001100100010;
            14'h431f: o_data_a = 16'b1110110000010000;
            14'h4320: o_data_a = 16'b0000000001011111;
            14'h4321: o_data_a = 16'b1110101010000111;
            14'h4322: o_data_a = 16'b0000000000000000;
            14'h4323: o_data_a = 16'b1111110010101000;
            14'h4324: o_data_a = 16'b1111110000010000;
            14'h4325: o_data_a = 16'b0000000000000101;
            14'h4326: o_data_a = 16'b1110001100001000;
            14'h4327: o_data_a = 16'b0000000001110111;
            14'h4328: o_data_a = 16'b1110110000010000;
            14'h4329: o_data_a = 16'b0000000000000000;
            14'h432a: o_data_a = 16'b1111110111101000;
            14'h432b: o_data_a = 16'b1110110010100000;
            14'h432c: o_data_a = 16'b1110001100001000;
            14'h432d: o_data_a = 16'b0000000000000000;
            14'h432e: o_data_a = 16'b1111110111001000;
            14'h432f: o_data_a = 16'b1111110010100000;
            14'h4330: o_data_a = 16'b1110101010001000;
            14'h4331: o_data_a = 16'b0000000000000000;
            14'h4332: o_data_a = 16'b1111110111001000;
            14'h4333: o_data_a = 16'b1111110010100000;
            14'h4334: o_data_a = 16'b1110101010001000;
            14'h4335: o_data_a = 16'b0000000000000000;
            14'h4336: o_data_a = 16'b1111110111001000;
            14'h4337: o_data_a = 16'b1111110010100000;
            14'h4338: o_data_a = 16'b1110101010001000;
            14'h4339: o_data_a = 16'b0000000000110011;
            14'h433a: o_data_a = 16'b1110110000010000;
            14'h433b: o_data_a = 16'b0000000000000000;
            14'h433c: o_data_a = 16'b1111110111101000;
            14'h433d: o_data_a = 16'b1110110010100000;
            14'h433e: o_data_a = 16'b1110001100001000;
            14'h433f: o_data_a = 16'b0000000000110011;
            14'h4340: o_data_a = 16'b1110110000010000;
            14'h4341: o_data_a = 16'b0000000000000000;
            14'h4342: o_data_a = 16'b1111110111101000;
            14'h4343: o_data_a = 16'b1110110010100000;
            14'h4344: o_data_a = 16'b1110001100001000;
            14'h4345: o_data_a = 16'b0000000000110011;
            14'h4346: o_data_a = 16'b1110110000010000;
            14'h4347: o_data_a = 16'b0000000000000000;
            14'h4348: o_data_a = 16'b1111110111101000;
            14'h4349: o_data_a = 16'b1110110010100000;
            14'h434a: o_data_a = 16'b1110001100001000;
            14'h434b: o_data_a = 16'b0000000000111111;
            14'h434c: o_data_a = 16'b1110110000010000;
            14'h434d: o_data_a = 16'b0000000000000000;
            14'h434e: o_data_a = 16'b1111110111101000;
            14'h434f: o_data_a = 16'b1110110010100000;
            14'h4350: o_data_a = 16'b1110001100001000;
            14'h4351: o_data_a = 16'b0000000000111111;
            14'h4352: o_data_a = 16'b1110110000010000;
            14'h4353: o_data_a = 16'b0000000000000000;
            14'h4354: o_data_a = 16'b1111110111101000;
            14'h4355: o_data_a = 16'b1110110010100000;
            14'h4356: o_data_a = 16'b1110001100001000;
            14'h4357: o_data_a = 16'b0000000000010010;
            14'h4358: o_data_a = 16'b1110110000010000;
            14'h4359: o_data_a = 16'b0000000000000000;
            14'h435a: o_data_a = 16'b1111110111101000;
            14'h435b: o_data_a = 16'b1110110010100000;
            14'h435c: o_data_a = 16'b1110001100001000;
            14'h435d: o_data_a = 16'b0000000000000000;
            14'h435e: o_data_a = 16'b1111110111001000;
            14'h435f: o_data_a = 16'b1111110010100000;
            14'h4360: o_data_a = 16'b1110101010001000;
            14'h4361: o_data_a = 16'b0000000000000000;
            14'h4362: o_data_a = 16'b1111110111001000;
            14'h4363: o_data_a = 16'b1111110010100000;
            14'h4364: o_data_a = 16'b1110101010001000;
            14'h4365: o_data_a = 16'b0000000000001100;
            14'h4366: o_data_a = 16'b1110110000010000;
            14'h4367: o_data_a = 16'b0000000000001101;
            14'h4368: o_data_a = 16'b1110001100001000;
            14'h4369: o_data_a = 16'b0100010110110011;
            14'h436a: o_data_a = 16'b1110110000010000;
            14'h436b: o_data_a = 16'b0000000000001110;
            14'h436c: o_data_a = 16'b1110001100001000;
            14'h436d: o_data_a = 16'b0100001101110001;
            14'h436e: o_data_a = 16'b1110110000010000;
            14'h436f: o_data_a = 16'b0000000001011111;
            14'h4370: o_data_a = 16'b1110101010000111;
            14'h4371: o_data_a = 16'b0000000000000000;
            14'h4372: o_data_a = 16'b1111110010101000;
            14'h4373: o_data_a = 16'b1111110000010000;
            14'h4374: o_data_a = 16'b0000000000000101;
            14'h4375: o_data_a = 16'b1110001100001000;
            14'h4376: o_data_a = 16'b0000000001111000;
            14'h4377: o_data_a = 16'b1110110000010000;
            14'h4378: o_data_a = 16'b0000000000000000;
            14'h4379: o_data_a = 16'b1111110111101000;
            14'h437a: o_data_a = 16'b1110110010100000;
            14'h437b: o_data_a = 16'b1110001100001000;
            14'h437c: o_data_a = 16'b0000000000000000;
            14'h437d: o_data_a = 16'b1111110111001000;
            14'h437e: o_data_a = 16'b1111110010100000;
            14'h437f: o_data_a = 16'b1110101010001000;
            14'h4380: o_data_a = 16'b0000000000000000;
            14'h4381: o_data_a = 16'b1111110111001000;
            14'h4382: o_data_a = 16'b1111110010100000;
            14'h4383: o_data_a = 16'b1110101010001000;
            14'h4384: o_data_a = 16'b0000000000000000;
            14'h4385: o_data_a = 16'b1111110111001000;
            14'h4386: o_data_a = 16'b1111110010100000;
            14'h4387: o_data_a = 16'b1110101010001000;
            14'h4388: o_data_a = 16'b0000000000110011;
            14'h4389: o_data_a = 16'b1110110000010000;
            14'h438a: o_data_a = 16'b0000000000000000;
            14'h438b: o_data_a = 16'b1111110111101000;
            14'h438c: o_data_a = 16'b1110110010100000;
            14'h438d: o_data_a = 16'b1110001100001000;
            14'h438e: o_data_a = 16'b0000000000011110;
            14'h438f: o_data_a = 16'b1110110000010000;
            14'h4390: o_data_a = 16'b0000000000000000;
            14'h4391: o_data_a = 16'b1111110111101000;
            14'h4392: o_data_a = 16'b1110110010100000;
            14'h4393: o_data_a = 16'b1110001100001000;
            14'h4394: o_data_a = 16'b0000000000001100;
            14'h4395: o_data_a = 16'b1110110000010000;
            14'h4396: o_data_a = 16'b0000000000000000;
            14'h4397: o_data_a = 16'b1111110111101000;
            14'h4398: o_data_a = 16'b1110110010100000;
            14'h4399: o_data_a = 16'b1110001100001000;
            14'h439a: o_data_a = 16'b0000000000001100;
            14'h439b: o_data_a = 16'b1110110000010000;
            14'h439c: o_data_a = 16'b0000000000000000;
            14'h439d: o_data_a = 16'b1111110111101000;
            14'h439e: o_data_a = 16'b1110110010100000;
            14'h439f: o_data_a = 16'b1110001100001000;
            14'h43a0: o_data_a = 16'b0000000000011110;
            14'h43a1: o_data_a = 16'b1110110000010000;
            14'h43a2: o_data_a = 16'b0000000000000000;
            14'h43a3: o_data_a = 16'b1111110111101000;
            14'h43a4: o_data_a = 16'b1110110010100000;
            14'h43a5: o_data_a = 16'b1110001100001000;
            14'h43a6: o_data_a = 16'b0000000000110011;
            14'h43a7: o_data_a = 16'b1110110000010000;
            14'h43a8: o_data_a = 16'b0000000000000000;
            14'h43a9: o_data_a = 16'b1111110111101000;
            14'h43aa: o_data_a = 16'b1110110010100000;
            14'h43ab: o_data_a = 16'b1110001100001000;
            14'h43ac: o_data_a = 16'b0000000000000000;
            14'h43ad: o_data_a = 16'b1111110111001000;
            14'h43ae: o_data_a = 16'b1111110010100000;
            14'h43af: o_data_a = 16'b1110101010001000;
            14'h43b0: o_data_a = 16'b0000000000000000;
            14'h43b1: o_data_a = 16'b1111110111001000;
            14'h43b2: o_data_a = 16'b1111110010100000;
            14'h43b3: o_data_a = 16'b1110101010001000;
            14'h43b4: o_data_a = 16'b0000000000001100;
            14'h43b5: o_data_a = 16'b1110110000010000;
            14'h43b6: o_data_a = 16'b0000000000001101;
            14'h43b7: o_data_a = 16'b1110001100001000;
            14'h43b8: o_data_a = 16'b0100010110110011;
            14'h43b9: o_data_a = 16'b1110110000010000;
            14'h43ba: o_data_a = 16'b0000000000001110;
            14'h43bb: o_data_a = 16'b1110001100001000;
            14'h43bc: o_data_a = 16'b0100001111000000;
            14'h43bd: o_data_a = 16'b1110110000010000;
            14'h43be: o_data_a = 16'b0000000001011111;
            14'h43bf: o_data_a = 16'b1110101010000111;
            14'h43c0: o_data_a = 16'b0000000000000000;
            14'h43c1: o_data_a = 16'b1111110010101000;
            14'h43c2: o_data_a = 16'b1111110000010000;
            14'h43c3: o_data_a = 16'b0000000000000101;
            14'h43c4: o_data_a = 16'b1110001100001000;
            14'h43c5: o_data_a = 16'b0000000001111001;
            14'h43c6: o_data_a = 16'b1110110000010000;
            14'h43c7: o_data_a = 16'b0000000000000000;
            14'h43c8: o_data_a = 16'b1111110111101000;
            14'h43c9: o_data_a = 16'b1110110010100000;
            14'h43ca: o_data_a = 16'b1110001100001000;
            14'h43cb: o_data_a = 16'b0000000000000000;
            14'h43cc: o_data_a = 16'b1111110111001000;
            14'h43cd: o_data_a = 16'b1111110010100000;
            14'h43ce: o_data_a = 16'b1110101010001000;
            14'h43cf: o_data_a = 16'b0000000000000000;
            14'h43d0: o_data_a = 16'b1111110111001000;
            14'h43d1: o_data_a = 16'b1111110010100000;
            14'h43d2: o_data_a = 16'b1110101010001000;
            14'h43d3: o_data_a = 16'b0000000000000000;
            14'h43d4: o_data_a = 16'b1111110111001000;
            14'h43d5: o_data_a = 16'b1111110010100000;
            14'h43d6: o_data_a = 16'b1110101010001000;
            14'h43d7: o_data_a = 16'b0000000000110011;
            14'h43d8: o_data_a = 16'b1110110000010000;
            14'h43d9: o_data_a = 16'b0000000000000000;
            14'h43da: o_data_a = 16'b1111110111101000;
            14'h43db: o_data_a = 16'b1110110010100000;
            14'h43dc: o_data_a = 16'b1110001100001000;
            14'h43dd: o_data_a = 16'b0000000000110011;
            14'h43de: o_data_a = 16'b1110110000010000;
            14'h43df: o_data_a = 16'b0000000000000000;
            14'h43e0: o_data_a = 16'b1111110111101000;
            14'h43e1: o_data_a = 16'b1110110010100000;
            14'h43e2: o_data_a = 16'b1110001100001000;
            14'h43e3: o_data_a = 16'b0000000000110011;
            14'h43e4: o_data_a = 16'b1110110000010000;
            14'h43e5: o_data_a = 16'b0000000000000000;
            14'h43e6: o_data_a = 16'b1111110111101000;
            14'h43e7: o_data_a = 16'b1110110010100000;
            14'h43e8: o_data_a = 16'b1110001100001000;
            14'h43e9: o_data_a = 16'b0000000000111110;
            14'h43ea: o_data_a = 16'b1110110000010000;
            14'h43eb: o_data_a = 16'b0000000000000000;
            14'h43ec: o_data_a = 16'b1111110111101000;
            14'h43ed: o_data_a = 16'b1110110010100000;
            14'h43ee: o_data_a = 16'b1110001100001000;
            14'h43ef: o_data_a = 16'b0000000000110000;
            14'h43f0: o_data_a = 16'b1110110000010000;
            14'h43f1: o_data_a = 16'b0000000000000000;
            14'h43f2: o_data_a = 16'b1111110111101000;
            14'h43f3: o_data_a = 16'b1110110010100000;
            14'h43f4: o_data_a = 16'b1110001100001000;
            14'h43f5: o_data_a = 16'b0000000000011000;
            14'h43f6: o_data_a = 16'b1110110000010000;
            14'h43f7: o_data_a = 16'b0000000000000000;
            14'h43f8: o_data_a = 16'b1111110111101000;
            14'h43f9: o_data_a = 16'b1110110010100000;
            14'h43fa: o_data_a = 16'b1110001100001000;
            14'h43fb: o_data_a = 16'b0000000000001111;
            14'h43fc: o_data_a = 16'b1110110000010000;
            14'h43fd: o_data_a = 16'b0000000000000000;
            14'h43fe: o_data_a = 16'b1111110111101000;
            14'h43ff: o_data_a = 16'b1110110010100000;
            14'h4400: o_data_a = 16'b1110001100001000;
            14'h4401: o_data_a = 16'b0000000000000000;
            14'h4402: o_data_a = 16'b1111110111001000;
            14'h4403: o_data_a = 16'b1111110010100000;
            14'h4404: o_data_a = 16'b1110101010001000;
            14'h4405: o_data_a = 16'b0000000000001100;
            14'h4406: o_data_a = 16'b1110110000010000;
            14'h4407: o_data_a = 16'b0000000000001101;
            14'h4408: o_data_a = 16'b1110001100001000;
            14'h4409: o_data_a = 16'b0100010110110011;
            14'h440a: o_data_a = 16'b1110110000010000;
            14'h440b: o_data_a = 16'b0000000000001110;
            14'h440c: o_data_a = 16'b1110001100001000;
            14'h440d: o_data_a = 16'b0100010000010001;
            14'h440e: o_data_a = 16'b1110110000010000;
            14'h440f: o_data_a = 16'b0000000001011111;
            14'h4410: o_data_a = 16'b1110101010000111;
            14'h4411: o_data_a = 16'b0000000000000000;
            14'h4412: o_data_a = 16'b1111110010101000;
            14'h4413: o_data_a = 16'b1111110000010000;
            14'h4414: o_data_a = 16'b0000000000000101;
            14'h4415: o_data_a = 16'b1110001100001000;
            14'h4416: o_data_a = 16'b0000000001111010;
            14'h4417: o_data_a = 16'b1110110000010000;
            14'h4418: o_data_a = 16'b0000000000000000;
            14'h4419: o_data_a = 16'b1111110111101000;
            14'h441a: o_data_a = 16'b1110110010100000;
            14'h441b: o_data_a = 16'b1110001100001000;
            14'h441c: o_data_a = 16'b0000000000000000;
            14'h441d: o_data_a = 16'b1111110111001000;
            14'h441e: o_data_a = 16'b1111110010100000;
            14'h441f: o_data_a = 16'b1110101010001000;
            14'h4420: o_data_a = 16'b0000000000000000;
            14'h4421: o_data_a = 16'b1111110111001000;
            14'h4422: o_data_a = 16'b1111110010100000;
            14'h4423: o_data_a = 16'b1110101010001000;
            14'h4424: o_data_a = 16'b0000000000000000;
            14'h4425: o_data_a = 16'b1111110111001000;
            14'h4426: o_data_a = 16'b1111110010100000;
            14'h4427: o_data_a = 16'b1110101010001000;
            14'h4428: o_data_a = 16'b0000000000111111;
            14'h4429: o_data_a = 16'b1110110000010000;
            14'h442a: o_data_a = 16'b0000000000000000;
            14'h442b: o_data_a = 16'b1111110111101000;
            14'h442c: o_data_a = 16'b1110110010100000;
            14'h442d: o_data_a = 16'b1110001100001000;
            14'h442e: o_data_a = 16'b0000000000011011;
            14'h442f: o_data_a = 16'b1110110000010000;
            14'h4430: o_data_a = 16'b0000000000000000;
            14'h4431: o_data_a = 16'b1111110111101000;
            14'h4432: o_data_a = 16'b1110110010100000;
            14'h4433: o_data_a = 16'b1110001100001000;
            14'h4434: o_data_a = 16'b0000000000001100;
            14'h4435: o_data_a = 16'b1110110000010000;
            14'h4436: o_data_a = 16'b0000000000000000;
            14'h4437: o_data_a = 16'b1111110111101000;
            14'h4438: o_data_a = 16'b1110110010100000;
            14'h4439: o_data_a = 16'b1110001100001000;
            14'h443a: o_data_a = 16'b0000000000000110;
            14'h443b: o_data_a = 16'b1110110000010000;
            14'h443c: o_data_a = 16'b0000000000000000;
            14'h443d: o_data_a = 16'b1111110111101000;
            14'h443e: o_data_a = 16'b1110110010100000;
            14'h443f: o_data_a = 16'b1110001100001000;
            14'h4440: o_data_a = 16'b0000000000110011;
            14'h4441: o_data_a = 16'b1110110000010000;
            14'h4442: o_data_a = 16'b0000000000000000;
            14'h4443: o_data_a = 16'b1111110111101000;
            14'h4444: o_data_a = 16'b1110110010100000;
            14'h4445: o_data_a = 16'b1110001100001000;
            14'h4446: o_data_a = 16'b0000000000111111;
            14'h4447: o_data_a = 16'b1110110000010000;
            14'h4448: o_data_a = 16'b0000000000000000;
            14'h4449: o_data_a = 16'b1111110111101000;
            14'h444a: o_data_a = 16'b1110110010100000;
            14'h444b: o_data_a = 16'b1110001100001000;
            14'h444c: o_data_a = 16'b0000000000000000;
            14'h444d: o_data_a = 16'b1111110111001000;
            14'h444e: o_data_a = 16'b1111110010100000;
            14'h444f: o_data_a = 16'b1110101010001000;
            14'h4450: o_data_a = 16'b0000000000000000;
            14'h4451: o_data_a = 16'b1111110111001000;
            14'h4452: o_data_a = 16'b1111110010100000;
            14'h4453: o_data_a = 16'b1110101010001000;
            14'h4454: o_data_a = 16'b0000000000001100;
            14'h4455: o_data_a = 16'b1110110000010000;
            14'h4456: o_data_a = 16'b0000000000001101;
            14'h4457: o_data_a = 16'b1110001100001000;
            14'h4458: o_data_a = 16'b0100010110110011;
            14'h4459: o_data_a = 16'b1110110000010000;
            14'h445a: o_data_a = 16'b0000000000001110;
            14'h445b: o_data_a = 16'b1110001100001000;
            14'h445c: o_data_a = 16'b0100010001100000;
            14'h445d: o_data_a = 16'b1110110000010000;
            14'h445e: o_data_a = 16'b0000000001011111;
            14'h445f: o_data_a = 16'b1110101010000111;
            14'h4460: o_data_a = 16'b0000000000000000;
            14'h4461: o_data_a = 16'b1111110010101000;
            14'h4462: o_data_a = 16'b1111110000010000;
            14'h4463: o_data_a = 16'b0000000000000101;
            14'h4464: o_data_a = 16'b1110001100001000;
            14'h4465: o_data_a = 16'b0000000001111011;
            14'h4466: o_data_a = 16'b1110110000010000;
            14'h4467: o_data_a = 16'b0000000000000000;
            14'h4468: o_data_a = 16'b1111110111101000;
            14'h4469: o_data_a = 16'b1110110010100000;
            14'h446a: o_data_a = 16'b1110001100001000;
            14'h446b: o_data_a = 16'b0000000000111000;
            14'h446c: o_data_a = 16'b1110110000010000;
            14'h446d: o_data_a = 16'b0000000000000000;
            14'h446e: o_data_a = 16'b1111110111101000;
            14'h446f: o_data_a = 16'b1110110010100000;
            14'h4470: o_data_a = 16'b1110001100001000;
            14'h4471: o_data_a = 16'b0000000000001100;
            14'h4472: o_data_a = 16'b1110110000010000;
            14'h4473: o_data_a = 16'b0000000000000000;
            14'h4474: o_data_a = 16'b1111110111101000;
            14'h4475: o_data_a = 16'b1110110010100000;
            14'h4476: o_data_a = 16'b1110001100001000;
            14'h4477: o_data_a = 16'b0000000000001100;
            14'h4478: o_data_a = 16'b1110110000010000;
            14'h4479: o_data_a = 16'b0000000000000000;
            14'h447a: o_data_a = 16'b1111110111101000;
            14'h447b: o_data_a = 16'b1110110010100000;
            14'h447c: o_data_a = 16'b1110001100001000;
            14'h447d: o_data_a = 16'b0000000000001100;
            14'h447e: o_data_a = 16'b1110110000010000;
            14'h447f: o_data_a = 16'b0000000000000000;
            14'h4480: o_data_a = 16'b1111110111101000;
            14'h4481: o_data_a = 16'b1110110010100000;
            14'h4482: o_data_a = 16'b1110001100001000;
            14'h4483: o_data_a = 16'b0000000000000111;
            14'h4484: o_data_a = 16'b1110110000010000;
            14'h4485: o_data_a = 16'b0000000000000000;
            14'h4486: o_data_a = 16'b1111110111101000;
            14'h4487: o_data_a = 16'b1110110010100000;
            14'h4488: o_data_a = 16'b1110001100001000;
            14'h4489: o_data_a = 16'b0000000000001100;
            14'h448a: o_data_a = 16'b1110110000010000;
            14'h448b: o_data_a = 16'b0000000000000000;
            14'h448c: o_data_a = 16'b1111110111101000;
            14'h448d: o_data_a = 16'b1110110010100000;
            14'h448e: o_data_a = 16'b1110001100001000;
            14'h448f: o_data_a = 16'b0000000000001100;
            14'h4490: o_data_a = 16'b1110110000010000;
            14'h4491: o_data_a = 16'b0000000000000000;
            14'h4492: o_data_a = 16'b1111110111101000;
            14'h4493: o_data_a = 16'b1110110010100000;
            14'h4494: o_data_a = 16'b1110001100001000;
            14'h4495: o_data_a = 16'b0000000000001100;
            14'h4496: o_data_a = 16'b1110110000010000;
            14'h4497: o_data_a = 16'b0000000000000000;
            14'h4498: o_data_a = 16'b1111110111101000;
            14'h4499: o_data_a = 16'b1110110010100000;
            14'h449a: o_data_a = 16'b1110001100001000;
            14'h449b: o_data_a = 16'b0000000000111000;
            14'h449c: o_data_a = 16'b1110110000010000;
            14'h449d: o_data_a = 16'b0000000000000000;
            14'h449e: o_data_a = 16'b1111110111101000;
            14'h449f: o_data_a = 16'b1110110010100000;
            14'h44a0: o_data_a = 16'b1110001100001000;
            14'h44a1: o_data_a = 16'b0000000000000000;
            14'h44a2: o_data_a = 16'b1111110111001000;
            14'h44a3: o_data_a = 16'b1111110010100000;
            14'h44a4: o_data_a = 16'b1110101010001000;
            14'h44a5: o_data_a = 16'b0000000000000000;
            14'h44a6: o_data_a = 16'b1111110111001000;
            14'h44a7: o_data_a = 16'b1111110010100000;
            14'h44a8: o_data_a = 16'b1110101010001000;
            14'h44a9: o_data_a = 16'b0000000000001100;
            14'h44aa: o_data_a = 16'b1110110000010000;
            14'h44ab: o_data_a = 16'b0000000000001101;
            14'h44ac: o_data_a = 16'b1110001100001000;
            14'h44ad: o_data_a = 16'b0100010110110011;
            14'h44ae: o_data_a = 16'b1110110000010000;
            14'h44af: o_data_a = 16'b0000000000001110;
            14'h44b0: o_data_a = 16'b1110001100001000;
            14'h44b1: o_data_a = 16'b0100010010110101;
            14'h44b2: o_data_a = 16'b1110110000010000;
            14'h44b3: o_data_a = 16'b0000000001011111;
            14'h44b4: o_data_a = 16'b1110101010000111;
            14'h44b5: o_data_a = 16'b0000000000000000;
            14'h44b6: o_data_a = 16'b1111110010101000;
            14'h44b7: o_data_a = 16'b1111110000010000;
            14'h44b8: o_data_a = 16'b0000000000000101;
            14'h44b9: o_data_a = 16'b1110001100001000;
            14'h44ba: o_data_a = 16'b0000000001111100;
            14'h44bb: o_data_a = 16'b1110110000010000;
            14'h44bc: o_data_a = 16'b0000000000000000;
            14'h44bd: o_data_a = 16'b1111110111101000;
            14'h44be: o_data_a = 16'b1110110010100000;
            14'h44bf: o_data_a = 16'b1110001100001000;
            14'h44c0: o_data_a = 16'b0000000000001100;
            14'h44c1: o_data_a = 16'b1110110000010000;
            14'h44c2: o_data_a = 16'b0000000000000000;
            14'h44c3: o_data_a = 16'b1111110111101000;
            14'h44c4: o_data_a = 16'b1110110010100000;
            14'h44c5: o_data_a = 16'b1110001100001000;
            14'h44c6: o_data_a = 16'b0000000000001100;
            14'h44c7: o_data_a = 16'b1110110000010000;
            14'h44c8: o_data_a = 16'b0000000000000000;
            14'h44c9: o_data_a = 16'b1111110111101000;
            14'h44ca: o_data_a = 16'b1110110010100000;
            14'h44cb: o_data_a = 16'b1110001100001000;
            14'h44cc: o_data_a = 16'b0000000000001100;
            14'h44cd: o_data_a = 16'b1110110000010000;
            14'h44ce: o_data_a = 16'b0000000000000000;
            14'h44cf: o_data_a = 16'b1111110111101000;
            14'h44d0: o_data_a = 16'b1110110010100000;
            14'h44d1: o_data_a = 16'b1110001100001000;
            14'h44d2: o_data_a = 16'b0000000000001100;
            14'h44d3: o_data_a = 16'b1110110000010000;
            14'h44d4: o_data_a = 16'b0000000000000000;
            14'h44d5: o_data_a = 16'b1111110111101000;
            14'h44d6: o_data_a = 16'b1110110010100000;
            14'h44d7: o_data_a = 16'b1110001100001000;
            14'h44d8: o_data_a = 16'b0000000000001100;
            14'h44d9: o_data_a = 16'b1110110000010000;
            14'h44da: o_data_a = 16'b0000000000000000;
            14'h44db: o_data_a = 16'b1111110111101000;
            14'h44dc: o_data_a = 16'b1110110010100000;
            14'h44dd: o_data_a = 16'b1110001100001000;
            14'h44de: o_data_a = 16'b0000000000001100;
            14'h44df: o_data_a = 16'b1110110000010000;
            14'h44e0: o_data_a = 16'b0000000000000000;
            14'h44e1: o_data_a = 16'b1111110111101000;
            14'h44e2: o_data_a = 16'b1110110010100000;
            14'h44e3: o_data_a = 16'b1110001100001000;
            14'h44e4: o_data_a = 16'b0000000000001100;
            14'h44e5: o_data_a = 16'b1110110000010000;
            14'h44e6: o_data_a = 16'b0000000000000000;
            14'h44e7: o_data_a = 16'b1111110111101000;
            14'h44e8: o_data_a = 16'b1110110010100000;
            14'h44e9: o_data_a = 16'b1110001100001000;
            14'h44ea: o_data_a = 16'b0000000000001100;
            14'h44eb: o_data_a = 16'b1110110000010000;
            14'h44ec: o_data_a = 16'b0000000000000000;
            14'h44ed: o_data_a = 16'b1111110111101000;
            14'h44ee: o_data_a = 16'b1110110010100000;
            14'h44ef: o_data_a = 16'b1110001100001000;
            14'h44f0: o_data_a = 16'b0000000000001100;
            14'h44f1: o_data_a = 16'b1110110000010000;
            14'h44f2: o_data_a = 16'b0000000000000000;
            14'h44f3: o_data_a = 16'b1111110111101000;
            14'h44f4: o_data_a = 16'b1110110010100000;
            14'h44f5: o_data_a = 16'b1110001100001000;
            14'h44f6: o_data_a = 16'b0000000000000000;
            14'h44f7: o_data_a = 16'b1111110111001000;
            14'h44f8: o_data_a = 16'b1111110010100000;
            14'h44f9: o_data_a = 16'b1110101010001000;
            14'h44fa: o_data_a = 16'b0000000000000000;
            14'h44fb: o_data_a = 16'b1111110111001000;
            14'h44fc: o_data_a = 16'b1111110010100000;
            14'h44fd: o_data_a = 16'b1110101010001000;
            14'h44fe: o_data_a = 16'b0000000000001100;
            14'h44ff: o_data_a = 16'b1110110000010000;
            14'h4500: o_data_a = 16'b0000000000001101;
            14'h4501: o_data_a = 16'b1110001100001000;
            14'h4502: o_data_a = 16'b0100010110110011;
            14'h4503: o_data_a = 16'b1110110000010000;
            14'h4504: o_data_a = 16'b0000000000001110;
            14'h4505: o_data_a = 16'b1110001100001000;
            14'h4506: o_data_a = 16'b0100010100001010;
            14'h4507: o_data_a = 16'b1110110000010000;
            14'h4508: o_data_a = 16'b0000000001011111;
            14'h4509: o_data_a = 16'b1110101010000111;
            14'h450a: o_data_a = 16'b0000000000000000;
            14'h450b: o_data_a = 16'b1111110010101000;
            14'h450c: o_data_a = 16'b1111110000010000;
            14'h450d: o_data_a = 16'b0000000000000101;
            14'h450e: o_data_a = 16'b1110001100001000;
            14'h450f: o_data_a = 16'b0000000001111101;
            14'h4510: o_data_a = 16'b1110110000010000;
            14'h4511: o_data_a = 16'b0000000000000000;
            14'h4512: o_data_a = 16'b1111110111101000;
            14'h4513: o_data_a = 16'b1110110010100000;
            14'h4514: o_data_a = 16'b1110001100001000;
            14'h4515: o_data_a = 16'b0000000000000111;
            14'h4516: o_data_a = 16'b1110110000010000;
            14'h4517: o_data_a = 16'b0000000000000000;
            14'h4518: o_data_a = 16'b1111110111101000;
            14'h4519: o_data_a = 16'b1110110010100000;
            14'h451a: o_data_a = 16'b1110001100001000;
            14'h451b: o_data_a = 16'b0000000000001100;
            14'h451c: o_data_a = 16'b1110110000010000;
            14'h451d: o_data_a = 16'b0000000000000000;
            14'h451e: o_data_a = 16'b1111110111101000;
            14'h451f: o_data_a = 16'b1110110010100000;
            14'h4520: o_data_a = 16'b1110001100001000;
            14'h4521: o_data_a = 16'b0000000000001100;
            14'h4522: o_data_a = 16'b1110110000010000;
            14'h4523: o_data_a = 16'b0000000000000000;
            14'h4524: o_data_a = 16'b1111110111101000;
            14'h4525: o_data_a = 16'b1110110010100000;
            14'h4526: o_data_a = 16'b1110001100001000;
            14'h4527: o_data_a = 16'b0000000000001100;
            14'h4528: o_data_a = 16'b1110110000010000;
            14'h4529: o_data_a = 16'b0000000000000000;
            14'h452a: o_data_a = 16'b1111110111101000;
            14'h452b: o_data_a = 16'b1110110010100000;
            14'h452c: o_data_a = 16'b1110001100001000;
            14'h452d: o_data_a = 16'b0000000000111000;
            14'h452e: o_data_a = 16'b1110110000010000;
            14'h452f: o_data_a = 16'b0000000000000000;
            14'h4530: o_data_a = 16'b1111110111101000;
            14'h4531: o_data_a = 16'b1110110010100000;
            14'h4532: o_data_a = 16'b1110001100001000;
            14'h4533: o_data_a = 16'b0000000000001100;
            14'h4534: o_data_a = 16'b1110110000010000;
            14'h4535: o_data_a = 16'b0000000000000000;
            14'h4536: o_data_a = 16'b1111110111101000;
            14'h4537: o_data_a = 16'b1110110010100000;
            14'h4538: o_data_a = 16'b1110001100001000;
            14'h4539: o_data_a = 16'b0000000000001100;
            14'h453a: o_data_a = 16'b1110110000010000;
            14'h453b: o_data_a = 16'b0000000000000000;
            14'h453c: o_data_a = 16'b1111110111101000;
            14'h453d: o_data_a = 16'b1110110010100000;
            14'h453e: o_data_a = 16'b1110001100001000;
            14'h453f: o_data_a = 16'b0000000000001100;
            14'h4540: o_data_a = 16'b1110110000010000;
            14'h4541: o_data_a = 16'b0000000000000000;
            14'h4542: o_data_a = 16'b1111110111101000;
            14'h4543: o_data_a = 16'b1110110010100000;
            14'h4544: o_data_a = 16'b1110001100001000;
            14'h4545: o_data_a = 16'b0000000000000111;
            14'h4546: o_data_a = 16'b1110110000010000;
            14'h4547: o_data_a = 16'b0000000000000000;
            14'h4548: o_data_a = 16'b1111110111101000;
            14'h4549: o_data_a = 16'b1110110010100000;
            14'h454a: o_data_a = 16'b1110001100001000;
            14'h454b: o_data_a = 16'b0000000000000000;
            14'h454c: o_data_a = 16'b1111110111001000;
            14'h454d: o_data_a = 16'b1111110010100000;
            14'h454e: o_data_a = 16'b1110101010001000;
            14'h454f: o_data_a = 16'b0000000000000000;
            14'h4550: o_data_a = 16'b1111110111001000;
            14'h4551: o_data_a = 16'b1111110010100000;
            14'h4552: o_data_a = 16'b1110101010001000;
            14'h4553: o_data_a = 16'b0000000000001100;
            14'h4554: o_data_a = 16'b1110110000010000;
            14'h4555: o_data_a = 16'b0000000000001101;
            14'h4556: o_data_a = 16'b1110001100001000;
            14'h4557: o_data_a = 16'b0100010110110011;
            14'h4558: o_data_a = 16'b1110110000010000;
            14'h4559: o_data_a = 16'b0000000000001110;
            14'h455a: o_data_a = 16'b1110001100001000;
            14'h455b: o_data_a = 16'b0100010101011111;
            14'h455c: o_data_a = 16'b1110110000010000;
            14'h455d: o_data_a = 16'b0000000001011111;
            14'h455e: o_data_a = 16'b1110101010000111;
            14'h455f: o_data_a = 16'b0000000000000000;
            14'h4560: o_data_a = 16'b1111110010101000;
            14'h4561: o_data_a = 16'b1111110000010000;
            14'h4562: o_data_a = 16'b0000000000000101;
            14'h4563: o_data_a = 16'b1110001100001000;
            14'h4564: o_data_a = 16'b0000000001111110;
            14'h4565: o_data_a = 16'b1110110000010000;
            14'h4566: o_data_a = 16'b0000000000000000;
            14'h4567: o_data_a = 16'b1111110111101000;
            14'h4568: o_data_a = 16'b1110110010100000;
            14'h4569: o_data_a = 16'b1110001100001000;
            14'h456a: o_data_a = 16'b0000000000100110;
            14'h456b: o_data_a = 16'b1110110000010000;
            14'h456c: o_data_a = 16'b0000000000000000;
            14'h456d: o_data_a = 16'b1111110111101000;
            14'h456e: o_data_a = 16'b1110110010100000;
            14'h456f: o_data_a = 16'b1110001100001000;
            14'h4570: o_data_a = 16'b0000000000101101;
            14'h4571: o_data_a = 16'b1110110000010000;
            14'h4572: o_data_a = 16'b0000000000000000;
            14'h4573: o_data_a = 16'b1111110111101000;
            14'h4574: o_data_a = 16'b1110110010100000;
            14'h4575: o_data_a = 16'b1110001100001000;
            14'h4576: o_data_a = 16'b0000000000011001;
            14'h4577: o_data_a = 16'b1110110000010000;
            14'h4578: o_data_a = 16'b0000000000000000;
            14'h4579: o_data_a = 16'b1111110111101000;
            14'h457a: o_data_a = 16'b1110110010100000;
            14'h457b: o_data_a = 16'b1110001100001000;
            14'h457c: o_data_a = 16'b0000000000000000;
            14'h457d: o_data_a = 16'b1111110111001000;
            14'h457e: o_data_a = 16'b1111110010100000;
            14'h457f: o_data_a = 16'b1110101010001000;
            14'h4580: o_data_a = 16'b0000000000000000;
            14'h4581: o_data_a = 16'b1111110111001000;
            14'h4582: o_data_a = 16'b1111110010100000;
            14'h4583: o_data_a = 16'b1110101010001000;
            14'h4584: o_data_a = 16'b0000000000000000;
            14'h4585: o_data_a = 16'b1111110111001000;
            14'h4586: o_data_a = 16'b1111110010100000;
            14'h4587: o_data_a = 16'b1110101010001000;
            14'h4588: o_data_a = 16'b0000000000000000;
            14'h4589: o_data_a = 16'b1111110111001000;
            14'h458a: o_data_a = 16'b1111110010100000;
            14'h458b: o_data_a = 16'b1110101010001000;
            14'h458c: o_data_a = 16'b0000000000000000;
            14'h458d: o_data_a = 16'b1111110111001000;
            14'h458e: o_data_a = 16'b1111110010100000;
            14'h458f: o_data_a = 16'b1110101010001000;
            14'h4590: o_data_a = 16'b0000000000000000;
            14'h4591: o_data_a = 16'b1111110111001000;
            14'h4592: o_data_a = 16'b1111110010100000;
            14'h4593: o_data_a = 16'b1110101010001000;
            14'h4594: o_data_a = 16'b0000000000000000;
            14'h4595: o_data_a = 16'b1111110111001000;
            14'h4596: o_data_a = 16'b1111110010100000;
            14'h4597: o_data_a = 16'b1110101010001000;
            14'h4598: o_data_a = 16'b0000000000000000;
            14'h4599: o_data_a = 16'b1111110111001000;
            14'h459a: o_data_a = 16'b1111110010100000;
            14'h459b: o_data_a = 16'b1110101010001000;
            14'h459c: o_data_a = 16'b0000000000001100;
            14'h459d: o_data_a = 16'b1110110000010000;
            14'h459e: o_data_a = 16'b0000000000001101;
            14'h459f: o_data_a = 16'b1110001100001000;
            14'h45a0: o_data_a = 16'b0100010110110011;
            14'h45a1: o_data_a = 16'b1110110000010000;
            14'h45a2: o_data_a = 16'b0000000000001110;
            14'h45a3: o_data_a = 16'b1110001100001000;
            14'h45a4: o_data_a = 16'b0100010110101000;
            14'h45a5: o_data_a = 16'b1110110000010000;
            14'h45a6: o_data_a = 16'b0000000001011111;
            14'h45a7: o_data_a = 16'b1110101010000111;
            14'h45a8: o_data_a = 16'b0000000000000000;
            14'h45a9: o_data_a = 16'b1111110010101000;
            14'h45aa: o_data_a = 16'b1111110000010000;
            14'h45ab: o_data_a = 16'b0000000000000101;
            14'h45ac: o_data_a = 16'b1110001100001000;
            14'h45ad: o_data_a = 16'b0000000000000000;
            14'h45ae: o_data_a = 16'b1111110111001000;
            14'h45af: o_data_a = 16'b1111110010100000;
            14'h45b0: o_data_a = 16'b1110101010001000;
            14'h45b1: o_data_a = 16'b0000000000110110;
            14'h45b2: o_data_a = 16'b1110101010000111;
            14'h45b3: o_data_a = 16'b0000000000000000;
            14'h45b4: o_data_a = 16'b1111110111101000;
            14'h45b5: o_data_a = 16'b1110110010100000;
            14'h45b6: o_data_a = 16'b1110101010001000;
            14'h45b7: o_data_a = 16'b0000000000001011;
            14'h45b8: o_data_a = 16'b1110110000010000;
            14'h45b9: o_data_a = 16'b0000000000000000;
            14'h45ba: o_data_a = 16'b1111110111101000;
            14'h45bb: o_data_a = 16'b1110110010100000;
            14'h45bc: o_data_a = 16'b1110001100001000;
            14'h45bd: o_data_a = 16'b0000000000000001;
            14'h45be: o_data_a = 16'b1110110000010000;
            14'h45bf: o_data_a = 16'b0000000000001101;
            14'h45c0: o_data_a = 16'b1110001100001000;
            14'h45c1: o_data_a = 16'b0001011010110000;
            14'h45c2: o_data_a = 16'b1110110000010000;
            14'h45c3: o_data_a = 16'b0000000000001110;
            14'h45c4: o_data_a = 16'b1110001100001000;
            14'h45c5: o_data_a = 16'b0100010111001001;
            14'h45c6: o_data_a = 16'b1110110000010000;
            14'h45c7: o_data_a = 16'b0000000001011111;
            14'h45c8: o_data_a = 16'b1110101010000111;
            14'h45c9: o_data_a = 16'b0000000000000000;
            14'h45ca: o_data_a = 16'b1111110010101000;
            14'h45cb: o_data_a = 16'b1111110000010000;
            14'h45cc: o_data_a = 16'b0000000000000001;
            14'h45cd: o_data_a = 16'b1111110000100000;
            14'h45ce: o_data_a = 16'b1110001100001000;
            14'h45cf: o_data_a = 16'b0000000000000010;
            14'h45d0: o_data_a = 16'b1111110000100000;
            14'h45d1: o_data_a = 16'b1111110000010000;
            14'h45d2: o_data_a = 16'b0000000000000000;
            14'h45d3: o_data_a = 16'b1111110111101000;
            14'h45d4: o_data_a = 16'b1110110010100000;
            14'h45d5: o_data_a = 16'b1110001100001000;
            14'h45d6: o_data_a = 16'b0000000000011001;
            14'h45d7: o_data_a = 16'b1111110000010000;
            14'h45d8: o_data_a = 16'b0000000000000000;
            14'h45d9: o_data_a = 16'b1111110111101000;
            14'h45da: o_data_a = 16'b1110110010100000;
            14'h45db: o_data_a = 16'b1110001100001000;
            14'h45dc: o_data_a = 16'b0000000000000000;
            14'h45dd: o_data_a = 16'b1111110010101000;
            14'h45de: o_data_a = 16'b1111110000010000;
            14'h45df: o_data_a = 16'b1110110010100000;
            14'h45e0: o_data_a = 16'b1111000010001000;
            14'h45e1: o_data_a = 16'b0000000000000001;
            14'h45e2: o_data_a = 16'b1111110000100000;
            14'h45e3: o_data_a = 16'b1111110000010000;
            14'h45e4: o_data_a = 16'b0000000000000000;
            14'h45e5: o_data_a = 16'b1111110111101000;
            14'h45e6: o_data_a = 16'b1110110010100000;
            14'h45e7: o_data_a = 16'b1110001100001000;
            14'h45e8: o_data_a = 16'b0000000000000000;
            14'h45e9: o_data_a = 16'b1111110010101000;
            14'h45ea: o_data_a = 16'b1111110000010000;
            14'h45eb: o_data_a = 16'b0000000000000101;
            14'h45ec: o_data_a = 16'b1110001100001000;
            14'h45ed: o_data_a = 16'b0000000000000000;
            14'h45ee: o_data_a = 16'b1111110010101000;
            14'h45ef: o_data_a = 16'b1111110000010000;
            14'h45f0: o_data_a = 16'b0000000000000100;
            14'h45f1: o_data_a = 16'b1110001100001000;
            14'h45f2: o_data_a = 16'b0000000000000101;
            14'h45f3: o_data_a = 16'b1111110000010000;
            14'h45f4: o_data_a = 16'b0000000000000000;
            14'h45f5: o_data_a = 16'b1111110111101000;
            14'h45f6: o_data_a = 16'b1110110010100000;
            14'h45f7: o_data_a = 16'b1110001100001000;
            14'h45f8: o_data_a = 16'b0000000000000000;
            14'h45f9: o_data_a = 16'b1111110010101000;
            14'h45fa: o_data_a = 16'b1111110000010000;
            14'h45fb: o_data_a = 16'b0000000000000100;
            14'h45fc: o_data_a = 16'b1111110000100000;
            14'h45fd: o_data_a = 16'b1110001100001000;
            14'h45fe: o_data_a = 16'b0000000000000000;
            14'h45ff: o_data_a = 16'b1111110111001000;
            14'h4600: o_data_a = 16'b1111110010100000;
            14'h4601: o_data_a = 16'b1110101010001000;
            14'h4602: o_data_a = 16'b0000000000000001;
            14'h4603: o_data_a = 16'b1111110000100000;
            14'h4604: o_data_a = 16'b1111110000010000;
            14'h4605: o_data_a = 16'b0000000000000000;
            14'h4606: o_data_a = 16'b1111110111101000;
            14'h4607: o_data_a = 16'b1110110010100000;
            14'h4608: o_data_a = 16'b1110001100001000;
            14'h4609: o_data_a = 16'b0000000000000000;
            14'h460a: o_data_a = 16'b1111110010101000;
            14'h460b: o_data_a = 16'b1111110000010000;
            14'h460c: o_data_a = 16'b1110110010100000;
            14'h460d: o_data_a = 16'b1111000010001000;
            14'h460e: o_data_a = 16'b0000000000000010;
            14'h460f: o_data_a = 16'b1111110111100000;
            14'h4610: o_data_a = 16'b1111110000010000;
            14'h4611: o_data_a = 16'b0000000000000000;
            14'h4612: o_data_a = 16'b1111110111101000;
            14'h4613: o_data_a = 16'b1110110010100000;
            14'h4614: o_data_a = 16'b1110001100001000;
            14'h4615: o_data_a = 16'b0000000000000000;
            14'h4616: o_data_a = 16'b1111110010101000;
            14'h4617: o_data_a = 16'b1111110000010000;
            14'h4618: o_data_a = 16'b0000000000000101;
            14'h4619: o_data_a = 16'b1110001100001000;
            14'h461a: o_data_a = 16'b0000000000000000;
            14'h461b: o_data_a = 16'b1111110010101000;
            14'h461c: o_data_a = 16'b1111110000010000;
            14'h461d: o_data_a = 16'b0000000000000100;
            14'h461e: o_data_a = 16'b1110001100001000;
            14'h461f: o_data_a = 16'b0000000000000101;
            14'h4620: o_data_a = 16'b1111110000010000;
            14'h4621: o_data_a = 16'b0000000000000000;
            14'h4622: o_data_a = 16'b1111110111101000;
            14'h4623: o_data_a = 16'b1110110010100000;
            14'h4624: o_data_a = 16'b1110001100001000;
            14'h4625: o_data_a = 16'b0000000000000000;
            14'h4626: o_data_a = 16'b1111110010101000;
            14'h4627: o_data_a = 16'b1111110000010000;
            14'h4628: o_data_a = 16'b0000000000000100;
            14'h4629: o_data_a = 16'b1111110000100000;
            14'h462a: o_data_a = 16'b1110001100001000;
            14'h462b: o_data_a = 16'b0000000000000000;
            14'h462c: o_data_a = 16'b1111110111001000;
            14'h462d: o_data_a = 16'b1111110010100000;
            14'h462e: o_data_a = 16'b1110111111001000;
            14'h462f: o_data_a = 16'b0000000000000001;
            14'h4630: o_data_a = 16'b1111110000100000;
            14'h4631: o_data_a = 16'b1111110000010000;
            14'h4632: o_data_a = 16'b0000000000000000;
            14'h4633: o_data_a = 16'b1111110111101000;
            14'h4634: o_data_a = 16'b1110110010100000;
            14'h4635: o_data_a = 16'b1110001100001000;
            14'h4636: o_data_a = 16'b0000000000000000;
            14'h4637: o_data_a = 16'b1111110010101000;
            14'h4638: o_data_a = 16'b1111110000010000;
            14'h4639: o_data_a = 16'b1110110010100000;
            14'h463a: o_data_a = 16'b1111000010001000;
            14'h463b: o_data_a = 16'b0000000000000010;
            14'h463c: o_data_a = 16'b1111110111100000;
            14'h463d: o_data_a = 16'b1110110111100000;
            14'h463e: o_data_a = 16'b1111110000010000;
            14'h463f: o_data_a = 16'b0000000000000000;
            14'h4640: o_data_a = 16'b1111110111101000;
            14'h4641: o_data_a = 16'b1110110010100000;
            14'h4642: o_data_a = 16'b1110001100001000;
            14'h4643: o_data_a = 16'b0000000000000000;
            14'h4644: o_data_a = 16'b1111110010101000;
            14'h4645: o_data_a = 16'b1111110000010000;
            14'h4646: o_data_a = 16'b0000000000000101;
            14'h4647: o_data_a = 16'b1110001100001000;
            14'h4648: o_data_a = 16'b0000000000000000;
            14'h4649: o_data_a = 16'b1111110010101000;
            14'h464a: o_data_a = 16'b1111110000010000;
            14'h464b: o_data_a = 16'b0000000000000100;
            14'h464c: o_data_a = 16'b1110001100001000;
            14'h464d: o_data_a = 16'b0000000000000101;
            14'h464e: o_data_a = 16'b1111110000010000;
            14'h464f: o_data_a = 16'b0000000000000000;
            14'h4650: o_data_a = 16'b1111110111101000;
            14'h4651: o_data_a = 16'b1110110010100000;
            14'h4652: o_data_a = 16'b1110001100001000;
            14'h4653: o_data_a = 16'b0000000000000000;
            14'h4654: o_data_a = 16'b1111110010101000;
            14'h4655: o_data_a = 16'b1111110000010000;
            14'h4656: o_data_a = 16'b0000000000000100;
            14'h4657: o_data_a = 16'b1111110000100000;
            14'h4658: o_data_a = 16'b1110001100001000;
            14'h4659: o_data_a = 16'b0000000000000010;
            14'h465a: o_data_a = 16'b1110110000010000;
            14'h465b: o_data_a = 16'b0000000000000000;
            14'h465c: o_data_a = 16'b1111110111101000;
            14'h465d: o_data_a = 16'b1110110010100000;
            14'h465e: o_data_a = 16'b1110001100001000;
            14'h465f: o_data_a = 16'b0000000000000001;
            14'h4660: o_data_a = 16'b1111110000100000;
            14'h4661: o_data_a = 16'b1111110000010000;
            14'h4662: o_data_a = 16'b0000000000000000;
            14'h4663: o_data_a = 16'b1111110111101000;
            14'h4664: o_data_a = 16'b1110110010100000;
            14'h4665: o_data_a = 16'b1110001100001000;
            14'h4666: o_data_a = 16'b0000000000000000;
            14'h4667: o_data_a = 16'b1111110010101000;
            14'h4668: o_data_a = 16'b1111110000010000;
            14'h4669: o_data_a = 16'b1110110010100000;
            14'h466a: o_data_a = 16'b1111000010001000;
            14'h466b: o_data_a = 16'b0000000000000010;
            14'h466c: o_data_a = 16'b1111110000010000;
            14'h466d: o_data_a = 16'b0000000000000011;
            14'h466e: o_data_a = 16'b1110000010100000;
            14'h466f: o_data_a = 16'b1111110000010000;
            14'h4670: o_data_a = 16'b0000000000000000;
            14'h4671: o_data_a = 16'b1111110111101000;
            14'h4672: o_data_a = 16'b1110110010100000;
            14'h4673: o_data_a = 16'b1110001100001000;
            14'h4674: o_data_a = 16'b0000000000000000;
            14'h4675: o_data_a = 16'b1111110010101000;
            14'h4676: o_data_a = 16'b1111110000010000;
            14'h4677: o_data_a = 16'b0000000000000101;
            14'h4678: o_data_a = 16'b1110001100001000;
            14'h4679: o_data_a = 16'b0000000000000000;
            14'h467a: o_data_a = 16'b1111110010101000;
            14'h467b: o_data_a = 16'b1111110000010000;
            14'h467c: o_data_a = 16'b0000000000000100;
            14'h467d: o_data_a = 16'b1110001100001000;
            14'h467e: o_data_a = 16'b0000000000000101;
            14'h467f: o_data_a = 16'b1111110000010000;
            14'h4680: o_data_a = 16'b0000000000000000;
            14'h4681: o_data_a = 16'b1111110111101000;
            14'h4682: o_data_a = 16'b1110110010100000;
            14'h4683: o_data_a = 16'b1110001100001000;
            14'h4684: o_data_a = 16'b0000000000000000;
            14'h4685: o_data_a = 16'b1111110010101000;
            14'h4686: o_data_a = 16'b1111110000010000;
            14'h4687: o_data_a = 16'b0000000000000100;
            14'h4688: o_data_a = 16'b1111110000100000;
            14'h4689: o_data_a = 16'b1110001100001000;
            14'h468a: o_data_a = 16'b0000000000000011;
            14'h468b: o_data_a = 16'b1110110000010000;
            14'h468c: o_data_a = 16'b0000000000000000;
            14'h468d: o_data_a = 16'b1111110111101000;
            14'h468e: o_data_a = 16'b1110110010100000;
            14'h468f: o_data_a = 16'b1110001100001000;
            14'h4690: o_data_a = 16'b0000000000000001;
            14'h4691: o_data_a = 16'b1111110000100000;
            14'h4692: o_data_a = 16'b1111110000010000;
            14'h4693: o_data_a = 16'b0000000000000000;
            14'h4694: o_data_a = 16'b1111110111101000;
            14'h4695: o_data_a = 16'b1110110010100000;
            14'h4696: o_data_a = 16'b1110001100001000;
            14'h4697: o_data_a = 16'b0000000000000000;
            14'h4698: o_data_a = 16'b1111110010101000;
            14'h4699: o_data_a = 16'b1111110000010000;
            14'h469a: o_data_a = 16'b1110110010100000;
            14'h469b: o_data_a = 16'b1111000010001000;
            14'h469c: o_data_a = 16'b0000000000000010;
            14'h469d: o_data_a = 16'b1111110000010000;
            14'h469e: o_data_a = 16'b0000000000000100;
            14'h469f: o_data_a = 16'b1110000010100000;
            14'h46a0: o_data_a = 16'b1111110000010000;
            14'h46a1: o_data_a = 16'b0000000000000000;
            14'h46a2: o_data_a = 16'b1111110111101000;
            14'h46a3: o_data_a = 16'b1110110010100000;
            14'h46a4: o_data_a = 16'b1110001100001000;
            14'h46a5: o_data_a = 16'b0000000000000000;
            14'h46a6: o_data_a = 16'b1111110010101000;
            14'h46a7: o_data_a = 16'b1111110000010000;
            14'h46a8: o_data_a = 16'b0000000000000101;
            14'h46a9: o_data_a = 16'b1110001100001000;
            14'h46aa: o_data_a = 16'b0000000000000000;
            14'h46ab: o_data_a = 16'b1111110010101000;
            14'h46ac: o_data_a = 16'b1111110000010000;
            14'h46ad: o_data_a = 16'b0000000000000100;
            14'h46ae: o_data_a = 16'b1110001100001000;
            14'h46af: o_data_a = 16'b0000000000000101;
            14'h46b0: o_data_a = 16'b1111110000010000;
            14'h46b1: o_data_a = 16'b0000000000000000;
            14'h46b2: o_data_a = 16'b1111110111101000;
            14'h46b3: o_data_a = 16'b1110110010100000;
            14'h46b4: o_data_a = 16'b1110001100001000;
            14'h46b5: o_data_a = 16'b0000000000000000;
            14'h46b6: o_data_a = 16'b1111110010101000;
            14'h46b7: o_data_a = 16'b1111110000010000;
            14'h46b8: o_data_a = 16'b0000000000000100;
            14'h46b9: o_data_a = 16'b1111110000100000;
            14'h46ba: o_data_a = 16'b1110001100001000;
            14'h46bb: o_data_a = 16'b0000000000000100;
            14'h46bc: o_data_a = 16'b1110110000010000;
            14'h46bd: o_data_a = 16'b0000000000000000;
            14'h46be: o_data_a = 16'b1111110111101000;
            14'h46bf: o_data_a = 16'b1110110010100000;
            14'h46c0: o_data_a = 16'b1110001100001000;
            14'h46c1: o_data_a = 16'b0000000000000001;
            14'h46c2: o_data_a = 16'b1111110000100000;
            14'h46c3: o_data_a = 16'b1111110000010000;
            14'h46c4: o_data_a = 16'b0000000000000000;
            14'h46c5: o_data_a = 16'b1111110111101000;
            14'h46c6: o_data_a = 16'b1110110010100000;
            14'h46c7: o_data_a = 16'b1110001100001000;
            14'h46c8: o_data_a = 16'b0000000000000000;
            14'h46c9: o_data_a = 16'b1111110010101000;
            14'h46ca: o_data_a = 16'b1111110000010000;
            14'h46cb: o_data_a = 16'b1110110010100000;
            14'h46cc: o_data_a = 16'b1111000010001000;
            14'h46cd: o_data_a = 16'b0000000000000010;
            14'h46ce: o_data_a = 16'b1111110000010000;
            14'h46cf: o_data_a = 16'b0000000000000101;
            14'h46d0: o_data_a = 16'b1110000010100000;
            14'h46d1: o_data_a = 16'b1111110000010000;
            14'h46d2: o_data_a = 16'b0000000000000000;
            14'h46d3: o_data_a = 16'b1111110111101000;
            14'h46d4: o_data_a = 16'b1110110010100000;
            14'h46d5: o_data_a = 16'b1110001100001000;
            14'h46d6: o_data_a = 16'b0000000000000000;
            14'h46d7: o_data_a = 16'b1111110010101000;
            14'h46d8: o_data_a = 16'b1111110000010000;
            14'h46d9: o_data_a = 16'b0000000000000101;
            14'h46da: o_data_a = 16'b1110001100001000;
            14'h46db: o_data_a = 16'b0000000000000000;
            14'h46dc: o_data_a = 16'b1111110010101000;
            14'h46dd: o_data_a = 16'b1111110000010000;
            14'h46de: o_data_a = 16'b0000000000000100;
            14'h46df: o_data_a = 16'b1110001100001000;
            14'h46e0: o_data_a = 16'b0000000000000101;
            14'h46e1: o_data_a = 16'b1111110000010000;
            14'h46e2: o_data_a = 16'b0000000000000000;
            14'h46e3: o_data_a = 16'b1111110111101000;
            14'h46e4: o_data_a = 16'b1110110010100000;
            14'h46e5: o_data_a = 16'b1110001100001000;
            14'h46e6: o_data_a = 16'b0000000000000000;
            14'h46e7: o_data_a = 16'b1111110010101000;
            14'h46e8: o_data_a = 16'b1111110000010000;
            14'h46e9: o_data_a = 16'b0000000000000100;
            14'h46ea: o_data_a = 16'b1111110000100000;
            14'h46eb: o_data_a = 16'b1110001100001000;
            14'h46ec: o_data_a = 16'b0000000000000101;
            14'h46ed: o_data_a = 16'b1110110000010000;
            14'h46ee: o_data_a = 16'b0000000000000000;
            14'h46ef: o_data_a = 16'b1111110111101000;
            14'h46f0: o_data_a = 16'b1110110010100000;
            14'h46f1: o_data_a = 16'b1110001100001000;
            14'h46f2: o_data_a = 16'b0000000000000001;
            14'h46f3: o_data_a = 16'b1111110000100000;
            14'h46f4: o_data_a = 16'b1111110000010000;
            14'h46f5: o_data_a = 16'b0000000000000000;
            14'h46f6: o_data_a = 16'b1111110111101000;
            14'h46f7: o_data_a = 16'b1110110010100000;
            14'h46f8: o_data_a = 16'b1110001100001000;
            14'h46f9: o_data_a = 16'b0000000000000000;
            14'h46fa: o_data_a = 16'b1111110010101000;
            14'h46fb: o_data_a = 16'b1111110000010000;
            14'h46fc: o_data_a = 16'b1110110010100000;
            14'h46fd: o_data_a = 16'b1111000010001000;
            14'h46fe: o_data_a = 16'b0000000000000010;
            14'h46ff: o_data_a = 16'b1111110000010000;
            14'h4700: o_data_a = 16'b0000000000000110;
            14'h4701: o_data_a = 16'b1110000010100000;
            14'h4702: o_data_a = 16'b1111110000010000;
            14'h4703: o_data_a = 16'b0000000000000000;
            14'h4704: o_data_a = 16'b1111110111101000;
            14'h4705: o_data_a = 16'b1110110010100000;
            14'h4706: o_data_a = 16'b1110001100001000;
            14'h4707: o_data_a = 16'b0000000000000000;
            14'h4708: o_data_a = 16'b1111110010101000;
            14'h4709: o_data_a = 16'b1111110000010000;
            14'h470a: o_data_a = 16'b0000000000000101;
            14'h470b: o_data_a = 16'b1110001100001000;
            14'h470c: o_data_a = 16'b0000000000000000;
            14'h470d: o_data_a = 16'b1111110010101000;
            14'h470e: o_data_a = 16'b1111110000010000;
            14'h470f: o_data_a = 16'b0000000000000100;
            14'h4710: o_data_a = 16'b1110001100001000;
            14'h4711: o_data_a = 16'b0000000000000101;
            14'h4712: o_data_a = 16'b1111110000010000;
            14'h4713: o_data_a = 16'b0000000000000000;
            14'h4714: o_data_a = 16'b1111110111101000;
            14'h4715: o_data_a = 16'b1110110010100000;
            14'h4716: o_data_a = 16'b1110001100001000;
            14'h4717: o_data_a = 16'b0000000000000000;
            14'h4718: o_data_a = 16'b1111110010101000;
            14'h4719: o_data_a = 16'b1111110000010000;
            14'h471a: o_data_a = 16'b0000000000000100;
            14'h471b: o_data_a = 16'b1111110000100000;
            14'h471c: o_data_a = 16'b1110001100001000;
            14'h471d: o_data_a = 16'b0000000000000110;
            14'h471e: o_data_a = 16'b1110110000010000;
            14'h471f: o_data_a = 16'b0000000000000000;
            14'h4720: o_data_a = 16'b1111110111101000;
            14'h4721: o_data_a = 16'b1110110010100000;
            14'h4722: o_data_a = 16'b1110001100001000;
            14'h4723: o_data_a = 16'b0000000000000001;
            14'h4724: o_data_a = 16'b1111110000100000;
            14'h4725: o_data_a = 16'b1111110000010000;
            14'h4726: o_data_a = 16'b0000000000000000;
            14'h4727: o_data_a = 16'b1111110111101000;
            14'h4728: o_data_a = 16'b1110110010100000;
            14'h4729: o_data_a = 16'b1110001100001000;
            14'h472a: o_data_a = 16'b0000000000000000;
            14'h472b: o_data_a = 16'b1111110010101000;
            14'h472c: o_data_a = 16'b1111110000010000;
            14'h472d: o_data_a = 16'b1110110010100000;
            14'h472e: o_data_a = 16'b1111000010001000;
            14'h472f: o_data_a = 16'b0000000000000010;
            14'h4730: o_data_a = 16'b1111110000010000;
            14'h4731: o_data_a = 16'b0000000000000111;
            14'h4732: o_data_a = 16'b1110000010100000;
            14'h4733: o_data_a = 16'b1111110000010000;
            14'h4734: o_data_a = 16'b0000000000000000;
            14'h4735: o_data_a = 16'b1111110111101000;
            14'h4736: o_data_a = 16'b1110110010100000;
            14'h4737: o_data_a = 16'b1110001100001000;
            14'h4738: o_data_a = 16'b0000000000000000;
            14'h4739: o_data_a = 16'b1111110010101000;
            14'h473a: o_data_a = 16'b1111110000010000;
            14'h473b: o_data_a = 16'b0000000000000101;
            14'h473c: o_data_a = 16'b1110001100001000;
            14'h473d: o_data_a = 16'b0000000000000000;
            14'h473e: o_data_a = 16'b1111110010101000;
            14'h473f: o_data_a = 16'b1111110000010000;
            14'h4740: o_data_a = 16'b0000000000000100;
            14'h4741: o_data_a = 16'b1110001100001000;
            14'h4742: o_data_a = 16'b0000000000000101;
            14'h4743: o_data_a = 16'b1111110000010000;
            14'h4744: o_data_a = 16'b0000000000000000;
            14'h4745: o_data_a = 16'b1111110111101000;
            14'h4746: o_data_a = 16'b1110110010100000;
            14'h4747: o_data_a = 16'b1110001100001000;
            14'h4748: o_data_a = 16'b0000000000000000;
            14'h4749: o_data_a = 16'b1111110010101000;
            14'h474a: o_data_a = 16'b1111110000010000;
            14'h474b: o_data_a = 16'b0000000000000100;
            14'h474c: o_data_a = 16'b1111110000100000;
            14'h474d: o_data_a = 16'b1110001100001000;
            14'h474e: o_data_a = 16'b0000000000000111;
            14'h474f: o_data_a = 16'b1110110000010000;
            14'h4750: o_data_a = 16'b0000000000000000;
            14'h4751: o_data_a = 16'b1111110111101000;
            14'h4752: o_data_a = 16'b1110110010100000;
            14'h4753: o_data_a = 16'b1110001100001000;
            14'h4754: o_data_a = 16'b0000000000000001;
            14'h4755: o_data_a = 16'b1111110000100000;
            14'h4756: o_data_a = 16'b1111110000010000;
            14'h4757: o_data_a = 16'b0000000000000000;
            14'h4758: o_data_a = 16'b1111110111101000;
            14'h4759: o_data_a = 16'b1110110010100000;
            14'h475a: o_data_a = 16'b1110001100001000;
            14'h475b: o_data_a = 16'b0000000000000000;
            14'h475c: o_data_a = 16'b1111110010101000;
            14'h475d: o_data_a = 16'b1111110000010000;
            14'h475e: o_data_a = 16'b1110110010100000;
            14'h475f: o_data_a = 16'b1111000010001000;
            14'h4760: o_data_a = 16'b0000000000000010;
            14'h4761: o_data_a = 16'b1111110000010000;
            14'h4762: o_data_a = 16'b0000000000001000;
            14'h4763: o_data_a = 16'b1110000010100000;
            14'h4764: o_data_a = 16'b1111110000010000;
            14'h4765: o_data_a = 16'b0000000000000000;
            14'h4766: o_data_a = 16'b1111110111101000;
            14'h4767: o_data_a = 16'b1110110010100000;
            14'h4768: o_data_a = 16'b1110001100001000;
            14'h4769: o_data_a = 16'b0000000000000000;
            14'h476a: o_data_a = 16'b1111110010101000;
            14'h476b: o_data_a = 16'b1111110000010000;
            14'h476c: o_data_a = 16'b0000000000000101;
            14'h476d: o_data_a = 16'b1110001100001000;
            14'h476e: o_data_a = 16'b0000000000000000;
            14'h476f: o_data_a = 16'b1111110010101000;
            14'h4770: o_data_a = 16'b1111110000010000;
            14'h4771: o_data_a = 16'b0000000000000100;
            14'h4772: o_data_a = 16'b1110001100001000;
            14'h4773: o_data_a = 16'b0000000000000101;
            14'h4774: o_data_a = 16'b1111110000010000;
            14'h4775: o_data_a = 16'b0000000000000000;
            14'h4776: o_data_a = 16'b1111110111101000;
            14'h4777: o_data_a = 16'b1110110010100000;
            14'h4778: o_data_a = 16'b1110001100001000;
            14'h4779: o_data_a = 16'b0000000000000000;
            14'h477a: o_data_a = 16'b1111110010101000;
            14'h477b: o_data_a = 16'b1111110000010000;
            14'h477c: o_data_a = 16'b0000000000000100;
            14'h477d: o_data_a = 16'b1111110000100000;
            14'h477e: o_data_a = 16'b1110001100001000;
            14'h477f: o_data_a = 16'b0000000000001000;
            14'h4780: o_data_a = 16'b1110110000010000;
            14'h4781: o_data_a = 16'b0000000000000000;
            14'h4782: o_data_a = 16'b1111110111101000;
            14'h4783: o_data_a = 16'b1110110010100000;
            14'h4784: o_data_a = 16'b1110001100001000;
            14'h4785: o_data_a = 16'b0000000000000001;
            14'h4786: o_data_a = 16'b1111110000100000;
            14'h4787: o_data_a = 16'b1111110000010000;
            14'h4788: o_data_a = 16'b0000000000000000;
            14'h4789: o_data_a = 16'b1111110111101000;
            14'h478a: o_data_a = 16'b1110110010100000;
            14'h478b: o_data_a = 16'b1110001100001000;
            14'h478c: o_data_a = 16'b0000000000000000;
            14'h478d: o_data_a = 16'b1111110010101000;
            14'h478e: o_data_a = 16'b1111110000010000;
            14'h478f: o_data_a = 16'b1110110010100000;
            14'h4790: o_data_a = 16'b1111000010001000;
            14'h4791: o_data_a = 16'b0000000000000010;
            14'h4792: o_data_a = 16'b1111110000010000;
            14'h4793: o_data_a = 16'b0000000000001001;
            14'h4794: o_data_a = 16'b1110000010100000;
            14'h4795: o_data_a = 16'b1111110000010000;
            14'h4796: o_data_a = 16'b0000000000000000;
            14'h4797: o_data_a = 16'b1111110111101000;
            14'h4798: o_data_a = 16'b1110110010100000;
            14'h4799: o_data_a = 16'b1110001100001000;
            14'h479a: o_data_a = 16'b0000000000000000;
            14'h479b: o_data_a = 16'b1111110010101000;
            14'h479c: o_data_a = 16'b1111110000010000;
            14'h479d: o_data_a = 16'b0000000000000101;
            14'h479e: o_data_a = 16'b1110001100001000;
            14'h479f: o_data_a = 16'b0000000000000000;
            14'h47a0: o_data_a = 16'b1111110010101000;
            14'h47a1: o_data_a = 16'b1111110000010000;
            14'h47a2: o_data_a = 16'b0000000000000100;
            14'h47a3: o_data_a = 16'b1110001100001000;
            14'h47a4: o_data_a = 16'b0000000000000101;
            14'h47a5: o_data_a = 16'b1111110000010000;
            14'h47a6: o_data_a = 16'b0000000000000000;
            14'h47a7: o_data_a = 16'b1111110111101000;
            14'h47a8: o_data_a = 16'b1110110010100000;
            14'h47a9: o_data_a = 16'b1110001100001000;
            14'h47aa: o_data_a = 16'b0000000000000000;
            14'h47ab: o_data_a = 16'b1111110010101000;
            14'h47ac: o_data_a = 16'b1111110000010000;
            14'h47ad: o_data_a = 16'b0000000000000100;
            14'h47ae: o_data_a = 16'b1111110000100000;
            14'h47af: o_data_a = 16'b1110001100001000;
            14'h47b0: o_data_a = 16'b0000000000001001;
            14'h47b1: o_data_a = 16'b1110110000010000;
            14'h47b2: o_data_a = 16'b0000000000000000;
            14'h47b3: o_data_a = 16'b1111110111101000;
            14'h47b4: o_data_a = 16'b1110110010100000;
            14'h47b5: o_data_a = 16'b1110001100001000;
            14'h47b6: o_data_a = 16'b0000000000000001;
            14'h47b7: o_data_a = 16'b1111110000100000;
            14'h47b8: o_data_a = 16'b1111110000010000;
            14'h47b9: o_data_a = 16'b0000000000000000;
            14'h47ba: o_data_a = 16'b1111110111101000;
            14'h47bb: o_data_a = 16'b1110110010100000;
            14'h47bc: o_data_a = 16'b1110001100001000;
            14'h47bd: o_data_a = 16'b0000000000000000;
            14'h47be: o_data_a = 16'b1111110010101000;
            14'h47bf: o_data_a = 16'b1111110000010000;
            14'h47c0: o_data_a = 16'b1110110010100000;
            14'h47c1: o_data_a = 16'b1111000010001000;
            14'h47c2: o_data_a = 16'b0000000000000010;
            14'h47c3: o_data_a = 16'b1111110000010000;
            14'h47c4: o_data_a = 16'b0000000000001010;
            14'h47c5: o_data_a = 16'b1110000010100000;
            14'h47c6: o_data_a = 16'b1111110000010000;
            14'h47c7: o_data_a = 16'b0000000000000000;
            14'h47c8: o_data_a = 16'b1111110111101000;
            14'h47c9: o_data_a = 16'b1110110010100000;
            14'h47ca: o_data_a = 16'b1110001100001000;
            14'h47cb: o_data_a = 16'b0000000000000000;
            14'h47cc: o_data_a = 16'b1111110010101000;
            14'h47cd: o_data_a = 16'b1111110000010000;
            14'h47ce: o_data_a = 16'b0000000000000101;
            14'h47cf: o_data_a = 16'b1110001100001000;
            14'h47d0: o_data_a = 16'b0000000000000000;
            14'h47d1: o_data_a = 16'b1111110010101000;
            14'h47d2: o_data_a = 16'b1111110000010000;
            14'h47d3: o_data_a = 16'b0000000000000100;
            14'h47d4: o_data_a = 16'b1110001100001000;
            14'h47d5: o_data_a = 16'b0000000000000101;
            14'h47d6: o_data_a = 16'b1111110000010000;
            14'h47d7: o_data_a = 16'b0000000000000000;
            14'h47d8: o_data_a = 16'b1111110111101000;
            14'h47d9: o_data_a = 16'b1110110010100000;
            14'h47da: o_data_a = 16'b1110001100001000;
            14'h47db: o_data_a = 16'b0000000000000000;
            14'h47dc: o_data_a = 16'b1111110010101000;
            14'h47dd: o_data_a = 16'b1111110000010000;
            14'h47de: o_data_a = 16'b0000000000000100;
            14'h47df: o_data_a = 16'b1111110000100000;
            14'h47e0: o_data_a = 16'b1110001100001000;
            14'h47e1: o_data_a = 16'b0000000000001010;
            14'h47e2: o_data_a = 16'b1110110000010000;
            14'h47e3: o_data_a = 16'b0000000000000000;
            14'h47e4: o_data_a = 16'b1111110111101000;
            14'h47e5: o_data_a = 16'b1110110010100000;
            14'h47e6: o_data_a = 16'b1110001100001000;
            14'h47e7: o_data_a = 16'b0000000000000001;
            14'h47e8: o_data_a = 16'b1111110000100000;
            14'h47e9: o_data_a = 16'b1111110000010000;
            14'h47ea: o_data_a = 16'b0000000000000000;
            14'h47eb: o_data_a = 16'b1111110111101000;
            14'h47ec: o_data_a = 16'b1110110010100000;
            14'h47ed: o_data_a = 16'b1110001100001000;
            14'h47ee: o_data_a = 16'b0000000000000000;
            14'h47ef: o_data_a = 16'b1111110010101000;
            14'h47f0: o_data_a = 16'b1111110000010000;
            14'h47f1: o_data_a = 16'b1110110010100000;
            14'h47f2: o_data_a = 16'b1111000010001000;
            14'h47f3: o_data_a = 16'b0000000000000010;
            14'h47f4: o_data_a = 16'b1111110000010000;
            14'h47f5: o_data_a = 16'b0000000000001011;
            14'h47f6: o_data_a = 16'b1110000010100000;
            14'h47f7: o_data_a = 16'b1111110000010000;
            14'h47f8: o_data_a = 16'b0000000000000000;
            14'h47f9: o_data_a = 16'b1111110111101000;
            14'h47fa: o_data_a = 16'b1110110010100000;
            14'h47fb: o_data_a = 16'b1110001100001000;
            14'h47fc: o_data_a = 16'b0000000000000000;
            14'h47fd: o_data_a = 16'b1111110010101000;
            14'h47fe: o_data_a = 16'b1111110000010000;
            14'h47ff: o_data_a = 16'b0000000000000101;
            14'h4800: o_data_a = 16'b1110001100001000;
            14'h4801: o_data_a = 16'b0000000000000000;
            14'h4802: o_data_a = 16'b1111110010101000;
            14'h4803: o_data_a = 16'b1111110000010000;
            14'h4804: o_data_a = 16'b0000000000000100;
            14'h4805: o_data_a = 16'b1110001100001000;
            14'h4806: o_data_a = 16'b0000000000000101;
            14'h4807: o_data_a = 16'b1111110000010000;
            14'h4808: o_data_a = 16'b0000000000000000;
            14'h4809: o_data_a = 16'b1111110111101000;
            14'h480a: o_data_a = 16'b1110110010100000;
            14'h480b: o_data_a = 16'b1110001100001000;
            14'h480c: o_data_a = 16'b0000000000000000;
            14'h480d: o_data_a = 16'b1111110010101000;
            14'h480e: o_data_a = 16'b1111110000010000;
            14'h480f: o_data_a = 16'b0000000000000100;
            14'h4810: o_data_a = 16'b1111110000100000;
            14'h4811: o_data_a = 16'b1110001100001000;
            14'h4812: o_data_a = 16'b0000000000000000;
            14'h4813: o_data_a = 16'b1111110111001000;
            14'h4814: o_data_a = 16'b1111110010100000;
            14'h4815: o_data_a = 16'b1110101010001000;
            14'h4816: o_data_a = 16'b0000000000110110;
            14'h4817: o_data_a = 16'b1110101010000111;
            14'h4818: o_data_a = 16'b0000000000000100;
            14'h4819: o_data_a = 16'b1110110000010000;
            14'h481a: o_data_a = 16'b1110001110010000;
            14'h481b: o_data_a = 16'b0000000000000000;
            14'h481c: o_data_a = 16'b1111110111101000;
            14'h481d: o_data_a = 16'b1110110010100000;
            14'h481e: o_data_a = 16'b1110101010001000;
            14'h481f: o_data_a = 16'b0100100000011010;
            14'h4820: o_data_a = 16'b1110001100000001;
            14'h4821: o_data_a = 16'b0000000001111111;
            14'h4822: o_data_a = 16'b1110110000010000;
            14'h4823: o_data_a = 16'b0000000000000000;
            14'h4824: o_data_a = 16'b1111110111101000;
            14'h4825: o_data_a = 16'b1110110010100000;
            14'h4826: o_data_a = 16'b1110001100001000;
            14'h4827: o_data_a = 16'b0000000000000001;
            14'h4828: o_data_a = 16'b1110110000010000;
            14'h4829: o_data_a = 16'b0000000000001101;
            14'h482a: o_data_a = 16'b1110001100001000;
            14'h482b: o_data_a = 16'b0001011010110000;
            14'h482c: o_data_a = 16'b1110110000010000;
            14'h482d: o_data_a = 16'b0000000000001110;
            14'h482e: o_data_a = 16'b1110001100001000;
            14'h482f: o_data_a = 16'b0100100000110011;
            14'h4830: o_data_a = 16'b1110110000010000;
            14'h4831: o_data_a = 16'b0000000001011111;
            14'h4832: o_data_a = 16'b1110101010000111;
            14'h4833: o_data_a = 16'b0000000000000000;
            14'h4834: o_data_a = 16'b1111110010101000;
            14'h4835: o_data_a = 16'b1111110000010000;
            14'h4836: o_data_a = 16'b0000000000011010;
            14'h4837: o_data_a = 16'b1110001100001000;
            14'h4838: o_data_a = 16'b0000000000000000;
            14'h4839: o_data_a = 16'b1111110111001000;
            14'h483a: o_data_a = 16'b1111110010100000;
            14'h483b: o_data_a = 16'b1110101010001000;
            14'h483c: o_data_a = 16'b0000000000000000;
            14'h483d: o_data_a = 16'b1111110010101000;
            14'h483e: o_data_a = 16'b1111110000010000;
            14'h483f: o_data_a = 16'b0000000000000001;
            14'h4840: o_data_a = 16'b1111110111100000;
            14'h4841: o_data_a = 16'b1110110111100000;
            14'h4842: o_data_a = 16'b1110001100001000;
            14'h4843: o_data_a = 16'b0000000000000001;
            14'h4844: o_data_a = 16'b1111110111100000;
            14'h4845: o_data_a = 16'b1110110111100000;
            14'h4846: o_data_a = 16'b1111110000010000;
            14'h4847: o_data_a = 16'b0000000000000000;
            14'h4848: o_data_a = 16'b1111110111101000;
            14'h4849: o_data_a = 16'b1110110010100000;
            14'h484a: o_data_a = 16'b1110001100001000;
            14'h484b: o_data_a = 16'b0000000001111111;
            14'h484c: o_data_a = 16'b1110110000010000;
            14'h484d: o_data_a = 16'b0000000000000000;
            14'h484e: o_data_a = 16'b1111110111101000;
            14'h484f: o_data_a = 16'b1110110010100000;
            14'h4850: o_data_a = 16'b1110001100001000;
            14'h4851: o_data_a = 16'b0100100001010101;
            14'h4852: o_data_a = 16'b1110110000010000;
            14'h4853: o_data_a = 16'b0000000000100110;
            14'h4854: o_data_a = 16'b1110101010000111;
            14'h4855: o_data_a = 16'b0000000000000000;
            14'h4856: o_data_a = 16'b1111110010100000;
            14'h4857: o_data_a = 16'b1111110001001000;
            14'h4858: o_data_a = 16'b0000000000000000;
            14'h4859: o_data_a = 16'b1111110010101000;
            14'h485a: o_data_a = 16'b1111110000010000;
            14'h485b: o_data_a = 16'b0100100110101011;
            14'h485c: o_data_a = 16'b1110001100000101;
            14'h485d: o_data_a = 16'b0000000000000001;
            14'h485e: o_data_a = 16'b1111110111100000;
            14'h485f: o_data_a = 16'b1110110111100000;
            14'h4860: o_data_a = 16'b1111110000010000;
            14'h4861: o_data_a = 16'b0000000000000000;
            14'h4862: o_data_a = 16'b1111110111101000;
            14'h4863: o_data_a = 16'b1110110010100000;
            14'h4864: o_data_a = 16'b1110001100001000;
            14'h4865: o_data_a = 16'b0000000000011001;
            14'h4866: o_data_a = 16'b1111110000010000;
            14'h4867: o_data_a = 16'b0000000000000000;
            14'h4868: o_data_a = 16'b1111110111101000;
            14'h4869: o_data_a = 16'b1110110010100000;
            14'h486a: o_data_a = 16'b1110001100001000;
            14'h486b: o_data_a = 16'b0000000000000000;
            14'h486c: o_data_a = 16'b1111110010101000;
            14'h486d: o_data_a = 16'b1111110000010000;
            14'h486e: o_data_a = 16'b1110110010100000;
            14'h486f: o_data_a = 16'b1111000010001000;
            14'h4870: o_data_a = 16'b0000000000000000;
            14'h4871: o_data_a = 16'b1111110010101000;
            14'h4872: o_data_a = 16'b1111110000010000;
            14'h4873: o_data_a = 16'b0000000000000100;
            14'h4874: o_data_a = 16'b1110001100001000;
            14'h4875: o_data_a = 16'b0000000000000100;
            14'h4876: o_data_a = 16'b1111110000100000;
            14'h4877: o_data_a = 16'b1111110000010000;
            14'h4878: o_data_a = 16'b0000000000000000;
            14'h4879: o_data_a = 16'b1111110111101000;
            14'h487a: o_data_a = 16'b1110110010100000;
            14'h487b: o_data_a = 16'b1110001100001000;
            14'h487c: o_data_a = 16'b0000000000000000;
            14'h487d: o_data_a = 16'b1111110010101000;
            14'h487e: o_data_a = 16'b1111110000010000;
            14'h487f: o_data_a = 16'b0000000000000001;
            14'h4880: o_data_a = 16'b1111110000100000;
            14'h4881: o_data_a = 16'b1110001100001000;
            14'h4882: o_data_a = 16'b0000000000001011;
            14'h4883: o_data_a = 16'b1110110000010000;
            14'h4884: o_data_a = 16'b0000000000000000;
            14'h4885: o_data_a = 16'b1111110111101000;
            14'h4886: o_data_a = 16'b1110110010100000;
            14'h4887: o_data_a = 16'b1110001100001000;
            14'h4888: o_data_a = 16'b0000000000000001;
            14'h4889: o_data_a = 16'b1110110000010000;
            14'h488a: o_data_a = 16'b0000000000001101;
            14'h488b: o_data_a = 16'b1110001100001000;
            14'h488c: o_data_a = 16'b0001011010110000;
            14'h488d: o_data_a = 16'b1110110000010000;
            14'h488e: o_data_a = 16'b0000000000001110;
            14'h488f: o_data_a = 16'b1110001100001000;
            14'h4890: o_data_a = 16'b0100100010010100;
            14'h4891: o_data_a = 16'b1110110000010000;
            14'h4892: o_data_a = 16'b0000000001011111;
            14'h4893: o_data_a = 16'b1110101010000111;
            14'h4894: o_data_a = 16'b0000000000000000;
            14'h4895: o_data_a = 16'b1111110010101000;
            14'h4896: o_data_a = 16'b1111110000010000;
            14'h4897: o_data_a = 16'b0000000000000001;
            14'h4898: o_data_a = 16'b1111110111100000;
            14'h4899: o_data_a = 16'b1110001100001000;
            14'h489a: o_data_a = 16'b0000000000000001;
            14'h489b: o_data_a = 16'b1111110111100000;
            14'h489c: o_data_a = 16'b1110110111100000;
            14'h489d: o_data_a = 16'b1111110000010000;
            14'h489e: o_data_a = 16'b0000000000000000;
            14'h489f: o_data_a = 16'b1111110111101000;
            14'h48a0: o_data_a = 16'b1110110010100000;
            14'h48a1: o_data_a = 16'b1110001100001000;
            14'h48a2: o_data_a = 16'b0000000000011010;
            14'h48a3: o_data_a = 16'b1111110000010000;
            14'h48a4: o_data_a = 16'b0000000000000000;
            14'h48a5: o_data_a = 16'b1111110111101000;
            14'h48a6: o_data_a = 16'b1110110010100000;
            14'h48a7: o_data_a = 16'b1110001100001000;
            14'h48a8: o_data_a = 16'b0000000000000000;
            14'h48a9: o_data_a = 16'b1111110010101000;
            14'h48aa: o_data_a = 16'b1111110000010000;
            14'h48ab: o_data_a = 16'b1110110010100000;
            14'h48ac: o_data_a = 16'b1111000010001000;
            14'h48ad: o_data_a = 16'b0000000000000001;
            14'h48ae: o_data_a = 16'b1111110111100000;
            14'h48af: o_data_a = 16'b1111110000010000;
            14'h48b0: o_data_a = 16'b0000000000000000;
            14'h48b1: o_data_a = 16'b1111110111101000;
            14'h48b2: o_data_a = 16'b1110110010100000;
            14'h48b3: o_data_a = 16'b1110001100001000;
            14'h48b4: o_data_a = 16'b0000000000000000;
            14'h48b5: o_data_a = 16'b1111110010101000;
            14'h48b6: o_data_a = 16'b1111110000010000;
            14'h48b7: o_data_a = 16'b0000000000000101;
            14'h48b8: o_data_a = 16'b1110001100001000;
            14'h48b9: o_data_a = 16'b0000000000000000;
            14'h48ba: o_data_a = 16'b1111110010101000;
            14'h48bb: o_data_a = 16'b1111110000010000;
            14'h48bc: o_data_a = 16'b0000000000000100;
            14'h48bd: o_data_a = 16'b1110001100001000;
            14'h48be: o_data_a = 16'b0000000000000101;
            14'h48bf: o_data_a = 16'b1111110000010000;
            14'h48c0: o_data_a = 16'b0000000000000000;
            14'h48c1: o_data_a = 16'b1111110111101000;
            14'h48c2: o_data_a = 16'b1110110010100000;
            14'h48c3: o_data_a = 16'b1110001100001000;
            14'h48c4: o_data_a = 16'b0000000000000000;
            14'h48c5: o_data_a = 16'b1111110010101000;
            14'h48c6: o_data_a = 16'b1111110000010000;
            14'h48c7: o_data_a = 16'b0000000000000100;
            14'h48c8: o_data_a = 16'b1111110000100000;
            14'h48c9: o_data_a = 16'b1110001100001000;
            14'h48ca: o_data_a = 16'b0000000000000000;
            14'h48cb: o_data_a = 16'b1111110111001000;
            14'h48cc: o_data_a = 16'b1111110010100000;
            14'h48cd: o_data_a = 16'b1110101010001000;
            14'h48ce: o_data_a = 16'b0000000000000000;
            14'h48cf: o_data_a = 16'b1111110010101000;
            14'h48d0: o_data_a = 16'b1111110000010000;
            14'h48d1: o_data_a = 16'b0000000000000001;
            14'h48d2: o_data_a = 16'b1111110111100000;
            14'h48d3: o_data_a = 16'b1110110111100000;
            14'h48d4: o_data_a = 16'b1110110111100000;
            14'h48d5: o_data_a = 16'b1110001100001000;
            14'h48d6: o_data_a = 16'b0000000000000001;
            14'h48d7: o_data_a = 16'b1111110000010000;
            14'h48d8: o_data_a = 16'b0000000000000011;
            14'h48d9: o_data_a = 16'b1110000010100000;
            14'h48da: o_data_a = 16'b1111110000010000;
            14'h48db: o_data_a = 16'b0000000000000000;
            14'h48dc: o_data_a = 16'b1111110111101000;
            14'h48dd: o_data_a = 16'b1110110010100000;
            14'h48de: o_data_a = 16'b1110001100001000;
            14'h48df: o_data_a = 16'b0000000000001011;
            14'h48e0: o_data_a = 16'b1110110000010000;
            14'h48e1: o_data_a = 16'b0000000000000000;
            14'h48e2: o_data_a = 16'b1111110111101000;
            14'h48e3: o_data_a = 16'b1110110010100000;
            14'h48e4: o_data_a = 16'b1110001100001000;
            14'h48e5: o_data_a = 16'b0100100011101001;
            14'h48e6: o_data_a = 16'b1110110000010000;
            14'h48e7: o_data_a = 16'b0000000000100110;
            14'h48e8: o_data_a = 16'b1110101010000111;
            14'h48e9: o_data_a = 16'b0000000000000000;
            14'h48ea: o_data_a = 16'b1111110010100000;
            14'h48eb: o_data_a = 16'b1111110001001000;
            14'h48ec: o_data_a = 16'b0000000000000000;
            14'h48ed: o_data_a = 16'b1111110010101000;
            14'h48ee: o_data_a = 16'b1111110000010000;
            14'h48ef: o_data_a = 16'b0100100101101011;
            14'h48f0: o_data_a = 16'b1110001100000101;
            14'h48f1: o_data_a = 16'b0000000000000001;
            14'h48f2: o_data_a = 16'b1111110000010000;
            14'h48f3: o_data_a = 16'b0000000000000011;
            14'h48f4: o_data_a = 16'b1110000010100000;
            14'h48f5: o_data_a = 16'b1111110000010000;
            14'h48f6: o_data_a = 16'b0000000000000000;
            14'h48f7: o_data_a = 16'b1111110111101000;
            14'h48f8: o_data_a = 16'b1110110010100000;
            14'h48f9: o_data_a = 16'b1110001100001000;
            14'h48fa: o_data_a = 16'b0000000000000001;
            14'h48fb: o_data_a = 16'b1111110111100000;
            14'h48fc: o_data_a = 16'b1111110000010000;
            14'h48fd: o_data_a = 16'b0000000000000000;
            14'h48fe: o_data_a = 16'b1111110111101000;
            14'h48ff: o_data_a = 16'b1110110010100000;
            14'h4900: o_data_a = 16'b1110001100001000;
            14'h4901: o_data_a = 16'b0000000000000000;
            14'h4902: o_data_a = 16'b1111110010101000;
            14'h4903: o_data_a = 16'b1111110000010000;
            14'h4904: o_data_a = 16'b1110110010100000;
            14'h4905: o_data_a = 16'b1111000010001000;
            14'h4906: o_data_a = 16'b0000000000000001;
            14'h4907: o_data_a = 16'b1111110000010000;
            14'h4908: o_data_a = 16'b0000000000000011;
            14'h4909: o_data_a = 16'b1110000010100000;
            14'h490a: o_data_a = 16'b1111110000010000;
            14'h490b: o_data_a = 16'b0000000000000000;
            14'h490c: o_data_a = 16'b1111110111101000;
            14'h490d: o_data_a = 16'b1110110010100000;
            14'h490e: o_data_a = 16'b1110001100001000;
            14'h490f: o_data_a = 16'b0000000000000001;
            14'h4910: o_data_a = 16'b1111110000100000;
            14'h4911: o_data_a = 16'b1111110000010000;
            14'h4912: o_data_a = 16'b0000000000000000;
            14'h4913: o_data_a = 16'b1111110111101000;
            14'h4914: o_data_a = 16'b1110110010100000;
            14'h4915: o_data_a = 16'b1110001100001000;
            14'h4916: o_data_a = 16'b0000000000000000;
            14'h4917: o_data_a = 16'b1111110010101000;
            14'h4918: o_data_a = 16'b1111110000010000;
            14'h4919: o_data_a = 16'b1110110010100000;
            14'h491a: o_data_a = 16'b1111000010001000;
            14'h491b: o_data_a = 16'b0000000000000000;
            14'h491c: o_data_a = 16'b1111110010101000;
            14'h491d: o_data_a = 16'b1111110000010000;
            14'h491e: o_data_a = 16'b0000000000000100;
            14'h491f: o_data_a = 16'b1110001100001000;
            14'h4920: o_data_a = 16'b0000000000000100;
            14'h4921: o_data_a = 16'b1111110000100000;
            14'h4922: o_data_a = 16'b1111110000010000;
            14'h4923: o_data_a = 16'b0000000000000000;
            14'h4924: o_data_a = 16'b1111110111101000;
            14'h4925: o_data_a = 16'b1110110010100000;
            14'h4926: o_data_a = 16'b1110001100001000;
            14'h4927: o_data_a = 16'b0000000100000000;
            14'h4928: o_data_a = 16'b1110110000010000;
            14'h4929: o_data_a = 16'b0000000000000000;
            14'h492a: o_data_a = 16'b1111110111101000;
            14'h492b: o_data_a = 16'b1110110010100000;
            14'h492c: o_data_a = 16'b1110001100001000;
            14'h492d: o_data_a = 16'b0000000000000010;
            14'h492e: o_data_a = 16'b1110110000010000;
            14'h492f: o_data_a = 16'b0000000000001101;
            14'h4930: o_data_a = 16'b1110001100001000;
            14'h4931: o_data_a = 16'b0001101010100110;
            14'h4932: o_data_a = 16'b1110110000010000;
            14'h4933: o_data_a = 16'b0000000000001110;
            14'h4934: o_data_a = 16'b1110001100001000;
            14'h4935: o_data_a = 16'b0100100100111001;
            14'h4936: o_data_a = 16'b1110110000010000;
            14'h4937: o_data_a = 16'b0000000001011111;
            14'h4938: o_data_a = 16'b1110101010000111;
            14'h4939: o_data_a = 16'b0000000000000000;
            14'h493a: o_data_a = 16'b1111110010101000;
            14'h493b: o_data_a = 16'b1111110000010000;
            14'h493c: o_data_a = 16'b0000000000000101;
            14'h493d: o_data_a = 16'b1110001100001000;
            14'h493e: o_data_a = 16'b0000000000000000;
            14'h493f: o_data_a = 16'b1111110010101000;
            14'h4940: o_data_a = 16'b1111110000010000;
            14'h4941: o_data_a = 16'b0000000000000100;
            14'h4942: o_data_a = 16'b1110001100001000;
            14'h4943: o_data_a = 16'b0000000000000101;
            14'h4944: o_data_a = 16'b1111110000010000;
            14'h4945: o_data_a = 16'b0000000000000000;
            14'h4946: o_data_a = 16'b1111110111101000;
            14'h4947: o_data_a = 16'b1110110010100000;
            14'h4948: o_data_a = 16'b1110001100001000;
            14'h4949: o_data_a = 16'b0000000000000000;
            14'h494a: o_data_a = 16'b1111110010101000;
            14'h494b: o_data_a = 16'b1111110000010000;
            14'h494c: o_data_a = 16'b0000000000000100;
            14'h494d: o_data_a = 16'b1111110000100000;
            14'h494e: o_data_a = 16'b1110001100001000;
            14'h494f: o_data_a = 16'b0000000000000001;
            14'h4950: o_data_a = 16'b1111110000010000;
            14'h4951: o_data_a = 16'b0000000000000011;
            14'h4952: o_data_a = 16'b1110000010100000;
            14'h4953: o_data_a = 16'b1111110000010000;
            14'h4954: o_data_a = 16'b0000000000000000;
            14'h4955: o_data_a = 16'b1111110111101000;
            14'h4956: o_data_a = 16'b1110110010100000;
            14'h4957: o_data_a = 16'b1110001100001000;
            14'h4958: o_data_a = 16'b0000000000000000;
            14'h4959: o_data_a = 16'b1111110111001000;
            14'h495a: o_data_a = 16'b1111110010100000;
            14'h495b: o_data_a = 16'b1110111111001000;
            14'h495c: o_data_a = 16'b0000000000000000;
            14'h495d: o_data_a = 16'b1111110010101000;
            14'h495e: o_data_a = 16'b1111110000010000;
            14'h495f: o_data_a = 16'b1110110010100000;
            14'h4960: o_data_a = 16'b1111000010001000;
            14'h4961: o_data_a = 16'b0000000000000000;
            14'h4962: o_data_a = 16'b1111110010101000;
            14'h4963: o_data_a = 16'b1111110000010000;
            14'h4964: o_data_a = 16'b0000000000000001;
            14'h4965: o_data_a = 16'b1111110111100000;
            14'h4966: o_data_a = 16'b1110110111100000;
            14'h4967: o_data_a = 16'b1110110111100000;
            14'h4968: o_data_a = 16'b1110001100001000;
            14'h4969: o_data_a = 16'b0100100011010110;
            14'h496a: o_data_a = 16'b1110101010000111;
            14'h496b: o_data_a = 16'b0000000000000001;
            14'h496c: o_data_a = 16'b1111110111100000;
            14'h496d: o_data_a = 16'b1110110111100000;
            14'h496e: o_data_a = 16'b1111110000010000;
            14'h496f: o_data_a = 16'b0000000000000000;
            14'h4970: o_data_a = 16'b1111110111101000;
            14'h4971: o_data_a = 16'b1110110010100000;
            14'h4972: o_data_a = 16'b1110001100001000;
            14'h4973: o_data_a = 16'b0000000000000000;
            14'h4974: o_data_a = 16'b1111110111001000;
            14'h4975: o_data_a = 16'b1111110010100000;
            14'h4976: o_data_a = 16'b1110101010001000;
            14'h4977: o_data_a = 16'b0100100101111011;
            14'h4978: o_data_a = 16'b1110110000010000;
            14'h4979: o_data_a = 16'b0000000000000110;
            14'h497a: o_data_a = 16'b1110101010000111;
            14'h497b: o_data_a = 16'b0000000000000000;
            14'h497c: o_data_a = 16'b1111110010101000;
            14'h497d: o_data_a = 16'b1111110000010000;
            14'h497e: o_data_a = 16'b0100100110000010;
            14'h497f: o_data_a = 16'b1110001100000101;
            14'h4980: o_data_a = 16'b0100100110010001;
            14'h4981: o_data_a = 16'b1110101010000111;
            14'h4982: o_data_a = 16'b0000000000100000;
            14'h4983: o_data_a = 16'b1110110000010000;
            14'h4984: o_data_a = 16'b0000000000000000;
            14'h4985: o_data_a = 16'b1111110111101000;
            14'h4986: o_data_a = 16'b1110110010100000;
            14'h4987: o_data_a = 16'b1110001100001000;
            14'h4988: o_data_a = 16'b0000000000000000;
            14'h4989: o_data_a = 16'b1111110010101000;
            14'h498a: o_data_a = 16'b1111110000010000;
            14'h498b: o_data_a = 16'b0000000000000001;
            14'h498c: o_data_a = 16'b1111110111100000;
            14'h498d: o_data_a = 16'b1110110111100000;
            14'h498e: o_data_a = 16'b1110001100001000;
            14'h498f: o_data_a = 16'b0100100110101001;
            14'h4990: o_data_a = 16'b1110101010000111;
            14'h4991: o_data_a = 16'b0000000000000001;
            14'h4992: o_data_a = 16'b1111110111100000;
            14'h4993: o_data_a = 16'b1110110111100000;
            14'h4994: o_data_a = 16'b1111110000010000;
            14'h4995: o_data_a = 16'b0000000000000000;
            14'h4996: o_data_a = 16'b1111110111101000;
            14'h4997: o_data_a = 16'b1110110010100000;
            14'h4998: o_data_a = 16'b1110001100001000;
            14'h4999: o_data_a = 16'b0000000000000000;
            14'h499a: o_data_a = 16'b1111110111001000;
            14'h499b: o_data_a = 16'b1111110010100000;
            14'h499c: o_data_a = 16'b1110111111001000;
            14'h499d: o_data_a = 16'b0000000000000000;
            14'h499e: o_data_a = 16'b1111110010101000;
            14'h499f: o_data_a = 16'b1111110000010000;
            14'h49a0: o_data_a = 16'b1110110010100000;
            14'h49a1: o_data_a = 16'b1111000010001000;
            14'h49a2: o_data_a = 16'b0000000000000000;
            14'h49a3: o_data_a = 16'b1111110010101000;
            14'h49a4: o_data_a = 16'b1111110000010000;
            14'h49a5: o_data_a = 16'b0000000000000001;
            14'h49a6: o_data_a = 16'b1111110111100000;
            14'h49a7: o_data_a = 16'b1110110111100000;
            14'h49a8: o_data_a = 16'b1110001100001000;
            14'h49a9: o_data_a = 16'b0100100001000011;
            14'h49aa: o_data_a = 16'b1110101010000111;
            14'h49ab: o_data_a = 16'b0000000000000000;
            14'h49ac: o_data_a = 16'b1111110111001000;
            14'h49ad: o_data_a = 16'b1111110010100000;
            14'h49ae: o_data_a = 16'b1110101010001000;
            14'h49af: o_data_a = 16'b0000000000110110;
            14'h49b0: o_data_a = 16'b1110101010000111;
            14'h49b1: o_data_a = 16'b0000000000000000;
            14'h49b2: o_data_a = 16'b1111110111101000;
            14'h49b3: o_data_a = 16'b1110110010100000;
            14'h49b4: o_data_a = 16'b1110101010001000;
            14'h49b5: o_data_a = 16'b0000000000000010;
            14'h49b6: o_data_a = 16'b1111110000100000;
            14'h49b7: o_data_a = 16'b1111110000010000;
            14'h49b8: o_data_a = 16'b0000000000000000;
            14'h49b9: o_data_a = 16'b1111110111101000;
            14'h49ba: o_data_a = 16'b1110110010100000;
            14'h49bb: o_data_a = 16'b1110001100001000;
            14'h49bc: o_data_a = 16'b0000000000100000;
            14'h49bd: o_data_a = 16'b1110110000010000;
            14'h49be: o_data_a = 16'b0000000000000000;
            14'h49bf: o_data_a = 16'b1111110111101000;
            14'h49c0: o_data_a = 16'b1110110010100000;
            14'h49c1: o_data_a = 16'b1110001100001000;
            14'h49c2: o_data_a = 16'b0100100111000110;
            14'h49c3: o_data_a = 16'b1110110000010000;
            14'h49c4: o_data_a = 16'b0000000000100110;
            14'h49c5: o_data_a = 16'b1110101010000111;
            14'h49c6: o_data_a = 16'b0000000000000010;
            14'h49c7: o_data_a = 16'b1111110000100000;
            14'h49c8: o_data_a = 16'b1111110000010000;
            14'h49c9: o_data_a = 16'b0000000000000000;
            14'h49ca: o_data_a = 16'b1111110111101000;
            14'h49cb: o_data_a = 16'b1110110010100000;
            14'h49cc: o_data_a = 16'b1110001100001000;
            14'h49cd: o_data_a = 16'b0000000001111110;
            14'h49ce: o_data_a = 16'b1110110000010000;
            14'h49cf: o_data_a = 16'b0000000000000000;
            14'h49d0: o_data_a = 16'b1111110111101000;
            14'h49d1: o_data_a = 16'b1110110010100000;
            14'h49d2: o_data_a = 16'b1110001100001000;
            14'h49d3: o_data_a = 16'b0100100111010111;
            14'h49d4: o_data_a = 16'b1110110000010000;
            14'h49d5: o_data_a = 16'b0000000000010110;
            14'h49d6: o_data_a = 16'b1110101010000111;
            14'h49d7: o_data_a = 16'b0000000000000000;
            14'h49d8: o_data_a = 16'b1111110010101000;
            14'h49d9: o_data_a = 16'b1111110000010000;
            14'h49da: o_data_a = 16'b1110110010100000;
            14'h49db: o_data_a = 16'b1111010101001000;
            14'h49dc: o_data_a = 16'b0000000000000000;
            14'h49dd: o_data_a = 16'b1111110010101000;
            14'h49de: o_data_a = 16'b1111110000010000;
            14'h49df: o_data_a = 16'b0100100111100011;
            14'h49e0: o_data_a = 16'b1110001100000101;
            14'h49e1: o_data_a = 16'b0100100111101101;
            14'h49e2: o_data_a = 16'b1110101010000111;
            14'h49e3: o_data_a = 16'b0000000000000000;
            14'h49e4: o_data_a = 16'b1111110111001000;
            14'h49e5: o_data_a = 16'b1111110010100000;
            14'h49e6: o_data_a = 16'b1110101010001000;
            14'h49e7: o_data_a = 16'b0000000000000000;
            14'h49e8: o_data_a = 16'b1111110010101000;
            14'h49e9: o_data_a = 16'b1111110000010000;
            14'h49ea: o_data_a = 16'b0000000000000010;
            14'h49eb: o_data_a = 16'b1111110000100000;
            14'h49ec: o_data_a = 16'b1110001100001000;
            14'h49ed: o_data_a = 16'b0000000000010101;
            14'h49ee: o_data_a = 16'b1111110000010000;
            14'h49ef: o_data_a = 16'b0000000000000000;
            14'h49f0: o_data_a = 16'b1111110111101000;
            14'h49f1: o_data_a = 16'b1110110010100000;
            14'h49f2: o_data_a = 16'b1110001100001000;
            14'h49f3: o_data_a = 16'b0000000000000000;
            14'h49f4: o_data_a = 16'b1111110010101000;
            14'h49f5: o_data_a = 16'b1111110000010000;
            14'h49f6: o_data_a = 16'b0100100111111010;
            14'h49f7: o_data_a = 16'b1110001100000101;
            14'h49f8: o_data_a = 16'b0100101000100000;
            14'h49f9: o_data_a = 16'b1110101010000111;
            14'h49fa: o_data_a = 16'b0000000000000010;
            14'h49fb: o_data_a = 16'b1111110000100000;
            14'h49fc: o_data_a = 16'b1111110000010000;
            14'h49fd: o_data_a = 16'b0000000000000000;
            14'h49fe: o_data_a = 16'b1111110111101000;
            14'h49ff: o_data_a = 16'b1110110010100000;
            14'h4a00: o_data_a = 16'b1110001100001000;
            14'h4a01: o_data_a = 16'b0000000000011001;
            14'h4a02: o_data_a = 16'b1111110000010000;
            14'h4a03: o_data_a = 16'b0000000000000000;
            14'h4a04: o_data_a = 16'b1111110111101000;
            14'h4a05: o_data_a = 16'b1110110010100000;
            14'h4a06: o_data_a = 16'b1110001100001000;
            14'h4a07: o_data_a = 16'b0000000000000000;
            14'h4a08: o_data_a = 16'b1111110010101000;
            14'h4a09: o_data_a = 16'b1111110000010000;
            14'h4a0a: o_data_a = 16'b1110110010100000;
            14'h4a0b: o_data_a = 16'b1111000010001000;
            14'h4a0c: o_data_a = 16'b0000000000000000;
            14'h4a0d: o_data_a = 16'b1111110010101000;
            14'h4a0e: o_data_a = 16'b1111110000010000;
            14'h4a0f: o_data_a = 16'b0000000000000100;
            14'h4a10: o_data_a = 16'b1110001100001000;
            14'h4a11: o_data_a = 16'b0000000000000100;
            14'h4a12: o_data_a = 16'b1111110000100000;
            14'h4a13: o_data_a = 16'b1111110000010000;
            14'h4a14: o_data_a = 16'b0000000000000000;
            14'h4a15: o_data_a = 16'b1111110111101000;
            14'h4a16: o_data_a = 16'b1110110010100000;
            14'h4a17: o_data_a = 16'b1110001100001000;
            14'h4a18: o_data_a = 16'b0000000000000000;
            14'h4a19: o_data_a = 16'b1111110010101000;
            14'h4a1a: o_data_a = 16'b1111110000010000;
            14'h4a1b: o_data_a = 16'b0000000000000001;
            14'h4a1c: o_data_a = 16'b1111110000100000;
            14'h4a1d: o_data_a = 16'b1110001100001000;
            14'h4a1e: o_data_a = 16'b0100101001000100;
            14'h4a1f: o_data_a = 16'b1110101010000111;
            14'h4a20: o_data_a = 16'b0000000000000010;
            14'h4a21: o_data_a = 16'b1111110000100000;
            14'h4a22: o_data_a = 16'b1111110000010000;
            14'h4a23: o_data_a = 16'b0000000000000000;
            14'h4a24: o_data_a = 16'b1111110111101000;
            14'h4a25: o_data_a = 16'b1110110010100000;
            14'h4a26: o_data_a = 16'b1110001100001000;
            14'h4a27: o_data_a = 16'b0000000000011010;
            14'h4a28: o_data_a = 16'b1111110000010000;
            14'h4a29: o_data_a = 16'b0000000000000000;
            14'h4a2a: o_data_a = 16'b1111110111101000;
            14'h4a2b: o_data_a = 16'b1110110010100000;
            14'h4a2c: o_data_a = 16'b1110001100001000;
            14'h4a2d: o_data_a = 16'b0000000000000000;
            14'h4a2e: o_data_a = 16'b1111110010101000;
            14'h4a2f: o_data_a = 16'b1111110000010000;
            14'h4a30: o_data_a = 16'b1110110010100000;
            14'h4a31: o_data_a = 16'b1111000010001000;
            14'h4a32: o_data_a = 16'b0000000000000000;
            14'h4a33: o_data_a = 16'b1111110010101000;
            14'h4a34: o_data_a = 16'b1111110000010000;
            14'h4a35: o_data_a = 16'b0000000000000100;
            14'h4a36: o_data_a = 16'b1110001100001000;
            14'h4a37: o_data_a = 16'b0000000000000100;
            14'h4a38: o_data_a = 16'b1111110000100000;
            14'h4a39: o_data_a = 16'b1111110000010000;
            14'h4a3a: o_data_a = 16'b0000000000000000;
            14'h4a3b: o_data_a = 16'b1111110111101000;
            14'h4a3c: o_data_a = 16'b1110110010100000;
            14'h4a3d: o_data_a = 16'b1110001100001000;
            14'h4a3e: o_data_a = 16'b0000000000000000;
            14'h4a3f: o_data_a = 16'b1111110010101000;
            14'h4a40: o_data_a = 16'b1111110000010000;
            14'h4a41: o_data_a = 16'b0000000000000001;
            14'h4a42: o_data_a = 16'b1111110000100000;
            14'h4a43: o_data_a = 16'b1110001100001000;
            14'h4a44: o_data_a = 16'b0000000000000001;
            14'h4a45: o_data_a = 16'b1111110000100000;
            14'h4a46: o_data_a = 16'b1111110000010000;
            14'h4a47: o_data_a = 16'b0000000000000000;
            14'h4a48: o_data_a = 16'b1111110111101000;
            14'h4a49: o_data_a = 16'b1110110010100000;
            14'h4a4a: o_data_a = 16'b1110001100001000;
            14'h4a4b: o_data_a = 16'b0000000000110110;
            14'h4a4c: o_data_a = 16'b1110101010000111;
            14'h4a4d: o_data_a = 16'b0000000000000100;
            14'h4a4e: o_data_a = 16'b1110110000010000;
            14'h4a4f: o_data_a = 16'b1110001110010000;
            14'h4a50: o_data_a = 16'b0000000000000000;
            14'h4a51: o_data_a = 16'b1111110111101000;
            14'h4a52: o_data_a = 16'b1110110010100000;
            14'h4a53: o_data_a = 16'b1110101010001000;
            14'h4a54: o_data_a = 16'b0100101001001111;
            14'h4a55: o_data_a = 16'b1110001100000001;
            14'h4a56: o_data_a = 16'b0000000000000010;
            14'h4a57: o_data_a = 16'b1111110000100000;
            14'h4a58: o_data_a = 16'b1111110000010000;
            14'h4a59: o_data_a = 16'b0000000000000000;
            14'h4a5a: o_data_a = 16'b1111110111101000;
            14'h4a5b: o_data_a = 16'b1110110010100000;
            14'h4a5c: o_data_a = 16'b1110001100001000;
            14'h4a5d: o_data_a = 16'b0000000000000001;
            14'h4a5e: o_data_a = 16'b1110110000010000;
            14'h4a5f: o_data_a = 16'b0000000000001101;
            14'h4a60: o_data_a = 16'b1110001100001000;
            14'h4a61: o_data_a = 16'b0100100110110001;
            14'h4a62: o_data_a = 16'b1110110000010000;
            14'h4a63: o_data_a = 16'b0000000000001110;
            14'h4a64: o_data_a = 16'b1110001100001000;
            14'h4a65: o_data_a = 16'b0100101001101001;
            14'h4a66: o_data_a = 16'b1110110000010000;
            14'h4a67: o_data_a = 16'b0000000001011111;
            14'h4a68: o_data_a = 16'b1110101010000111;
            14'h4a69: o_data_a = 16'b0000000000000000;
            14'h4a6a: o_data_a = 16'b1111110010101000;
            14'h4a6b: o_data_a = 16'b1111110000010000;
            14'h4a6c: o_data_a = 16'b0000000000000001;
            14'h4a6d: o_data_a = 16'b1111110111100000;
            14'h4a6e: o_data_a = 16'b1110110111100000;
            14'h4a6f: o_data_a = 16'b1110001100001000;
            14'h4a70: o_data_a = 16'b0000000000010110;
            14'h4a71: o_data_a = 16'b1111110000010000;
            14'h4a72: o_data_a = 16'b0000000000000000;
            14'h4a73: o_data_a = 16'b1111110111101000;
            14'h4a74: o_data_a = 16'b1110110010100000;
            14'h4a75: o_data_a = 16'b1110001100001000;
            14'h4a76: o_data_a = 16'b0000000000000000;
            14'h4a77: o_data_a = 16'b1111110010101000;
            14'h4a78: o_data_a = 16'b1111110000010000;
            14'h4a79: o_data_a = 16'b0000000000000001;
            14'h4a7a: o_data_a = 16'b1111110000100000;
            14'h4a7b: o_data_a = 16'b1110001100001000;
            14'h4a7c: o_data_a = 16'b0000000000000001;
            14'h4a7d: o_data_a = 16'b1111110111100000;
            14'h4a7e: o_data_a = 16'b1111110000010000;
            14'h4a7f: o_data_a = 16'b0000000000000000;
            14'h4a80: o_data_a = 16'b1111110111101000;
            14'h4a81: o_data_a = 16'b1110110010100000;
            14'h4a82: o_data_a = 16'b1110001100001000;
            14'h4a83: o_data_a = 16'b0000000000001011;
            14'h4a84: o_data_a = 16'b1110110000010000;
            14'h4a85: o_data_a = 16'b0000000000000000;
            14'h4a86: o_data_a = 16'b1111110111101000;
            14'h4a87: o_data_a = 16'b1110110010100000;
            14'h4a88: o_data_a = 16'b1110001100001000;
            14'h4a89: o_data_a = 16'b0100101010001101;
            14'h4a8a: o_data_a = 16'b1110110000010000;
            14'h4a8b: o_data_a = 16'b0000000000100110;
            14'h4a8c: o_data_a = 16'b1110101010000111;
            14'h4a8d: o_data_a = 16'b0000000000000000;
            14'h4a8e: o_data_a = 16'b1111110010100000;
            14'h4a8f: o_data_a = 16'b1111110001001000;
            14'h4a90: o_data_a = 16'b0000000000000000;
            14'h4a91: o_data_a = 16'b1111110010101000;
            14'h4a92: o_data_a = 16'b1111110000010000;
            14'h4a93: o_data_a = 16'b0100101110010000;
            14'h4a94: o_data_a = 16'b1110001100000101;
            14'h4a95: o_data_a = 16'b0000000000010101;
            14'h4a96: o_data_a = 16'b1111110000010000;
            14'h4a97: o_data_a = 16'b0000000000000000;
            14'h4a98: o_data_a = 16'b1111110111101000;
            14'h4a99: o_data_a = 16'b1110110010100000;
            14'h4a9a: o_data_a = 16'b1110001100001000;
            14'h4a9b: o_data_a = 16'b0000000000000000;
            14'h4a9c: o_data_a = 16'b1111110010101000;
            14'h4a9d: o_data_a = 16'b1111110000010000;
            14'h4a9e: o_data_a = 16'b0100101010100010;
            14'h4a9f: o_data_a = 16'b1110001100000101;
            14'h4aa0: o_data_a = 16'b0100101011011001;
            14'h4aa1: o_data_a = 16'b1110101010000111;
            14'h4aa2: o_data_a = 16'b0000000000000001;
            14'h4aa3: o_data_a = 16'b1111110000100000;
            14'h4aa4: o_data_a = 16'b1111110000010000;
            14'h4aa5: o_data_a = 16'b0000000000000000;
            14'h4aa6: o_data_a = 16'b1111110111101000;
            14'h4aa7: o_data_a = 16'b1110110010100000;
            14'h4aa8: o_data_a = 16'b1110001100001000;
            14'h4aa9: o_data_a = 16'b0000000000010100;
            14'h4aaa: o_data_a = 16'b1111110000010000;
            14'h4aab: o_data_a = 16'b0000000000000000;
            14'h4aac: o_data_a = 16'b1111110111101000;
            14'h4aad: o_data_a = 16'b1110110010100000;
            14'h4aae: o_data_a = 16'b1110001100001000;
            14'h4aaf: o_data_a = 16'b0000000000000000;
            14'h4ab0: o_data_a = 16'b1111110010101000;
            14'h4ab1: o_data_a = 16'b1111110000010000;
            14'h4ab2: o_data_a = 16'b1110110010100000;
            14'h4ab3: o_data_a = 16'b1111000010001000;
            14'h4ab4: o_data_a = 16'b0000000000000000;
            14'h4ab5: o_data_a = 16'b1111110010101000;
            14'h4ab6: o_data_a = 16'b1111110000010000;
            14'h4ab7: o_data_a = 16'b0000000000000100;
            14'h4ab8: o_data_a = 16'b1110001100001000;
            14'h4ab9: o_data_a = 16'b0000000000000100;
            14'h4aba: o_data_a = 16'b1111110000100000;
            14'h4abb: o_data_a = 16'b1111110000010000;
            14'h4abc: o_data_a = 16'b0000000000000000;
            14'h4abd: o_data_a = 16'b1111110111101000;
            14'h4abe: o_data_a = 16'b1110110010100000;
            14'h4abf: o_data_a = 16'b1110001100001000;
            14'h4ac0: o_data_a = 16'b0000000100000000;
            14'h4ac1: o_data_a = 16'b1110110000010000;
            14'h4ac2: o_data_a = 16'b0000000000000000;
            14'h4ac3: o_data_a = 16'b1111110111101000;
            14'h4ac4: o_data_a = 16'b1110110010100000;
            14'h4ac5: o_data_a = 16'b1110001100001000;
            14'h4ac6: o_data_a = 16'b0000000000000000;
            14'h4ac7: o_data_a = 16'b1111110010100000;
            14'h4ac8: o_data_a = 16'b1111110001010000;
            14'h4ac9: o_data_a = 16'b1110011111001000;
            14'h4aca: o_data_a = 16'b0000000000000000;
            14'h4acb: o_data_a = 16'b1111110010101000;
            14'h4acc: o_data_a = 16'b1111110000010000;
            14'h4acd: o_data_a = 16'b1110110010100000;
            14'h4ace: o_data_a = 16'b1111000000001000;
            14'h4acf: o_data_a = 16'b0000000000000000;
            14'h4ad0: o_data_a = 16'b1111110010101000;
            14'h4ad1: o_data_a = 16'b1111110000010000;
            14'h4ad2: o_data_a = 16'b0000000000000001;
            14'h4ad3: o_data_a = 16'b1111110111100000;
            14'h4ad4: o_data_a = 16'b1110110111100000;
            14'h4ad5: o_data_a = 16'b1110110111100000;
            14'h4ad6: o_data_a = 16'b1110001100001000;
            14'h4ad7: o_data_a = 16'b0100101100001010;
            14'h4ad8: o_data_a = 16'b1110101010000111;
            14'h4ad9: o_data_a = 16'b0000000000000001;
            14'h4ada: o_data_a = 16'b1111110000100000;
            14'h4adb: o_data_a = 16'b1111110000010000;
            14'h4adc: o_data_a = 16'b0000000000000000;
            14'h4add: o_data_a = 16'b1111110111101000;
            14'h4ade: o_data_a = 16'b1110110010100000;
            14'h4adf: o_data_a = 16'b1110001100001000;
            14'h4ae0: o_data_a = 16'b0000000000010100;
            14'h4ae1: o_data_a = 16'b1111110000010000;
            14'h4ae2: o_data_a = 16'b0000000000000000;
            14'h4ae3: o_data_a = 16'b1111110111101000;
            14'h4ae4: o_data_a = 16'b1110110010100000;
            14'h4ae5: o_data_a = 16'b1110001100001000;
            14'h4ae6: o_data_a = 16'b0000000000000000;
            14'h4ae7: o_data_a = 16'b1111110010101000;
            14'h4ae8: o_data_a = 16'b1111110000010000;
            14'h4ae9: o_data_a = 16'b1110110010100000;
            14'h4aea: o_data_a = 16'b1111000010001000;
            14'h4aeb: o_data_a = 16'b0000000000000000;
            14'h4aec: o_data_a = 16'b1111110010101000;
            14'h4aed: o_data_a = 16'b1111110000010000;
            14'h4aee: o_data_a = 16'b0000000000000100;
            14'h4aef: o_data_a = 16'b1110001100001000;
            14'h4af0: o_data_a = 16'b0000000000000100;
            14'h4af1: o_data_a = 16'b1111110000100000;
            14'h4af2: o_data_a = 16'b1111110000010000;
            14'h4af3: o_data_a = 16'b0000000000000000;
            14'h4af4: o_data_a = 16'b1111110111101000;
            14'h4af5: o_data_a = 16'b1110110010100000;
            14'h4af6: o_data_a = 16'b1110001100001000;
            14'h4af7: o_data_a = 16'b0000000011111111;
            14'h4af8: o_data_a = 16'b1110110000010000;
            14'h4af9: o_data_a = 16'b0000000000000000;
            14'h4afa: o_data_a = 16'b1111110111101000;
            14'h4afb: o_data_a = 16'b1110110010100000;
            14'h4afc: o_data_a = 16'b1110001100001000;
            14'h4afd: o_data_a = 16'b0000000000000000;
            14'h4afe: o_data_a = 16'b1111110010101000;
            14'h4aff: o_data_a = 16'b1111110000010000;
            14'h4b00: o_data_a = 16'b1110110010100000;
            14'h4b01: o_data_a = 16'b1111000000001000;
            14'h4b02: o_data_a = 16'b0000000000000000;
            14'h4b03: o_data_a = 16'b1111110010101000;
            14'h4b04: o_data_a = 16'b1111110000010000;
            14'h4b05: o_data_a = 16'b0000000000000001;
            14'h4b06: o_data_a = 16'b1111110111100000;
            14'h4b07: o_data_a = 16'b1110110111100000;
            14'h4b08: o_data_a = 16'b1110110111100000;
            14'h4b09: o_data_a = 16'b1110001100001000;
            14'h4b0a: o_data_a = 16'b0000000000000001;
            14'h4b0b: o_data_a = 16'b1111110000100000;
            14'h4b0c: o_data_a = 16'b1111110000010000;
            14'h4b0d: o_data_a = 16'b0000000000000000;
            14'h4b0e: o_data_a = 16'b1111110111101000;
            14'h4b0f: o_data_a = 16'b1110110010100000;
            14'h4b10: o_data_a = 16'b1110001100001000;
            14'h4b11: o_data_a = 16'b0000000000010100;
            14'h4b12: o_data_a = 16'b1111110000010000;
            14'h4b13: o_data_a = 16'b0000000000000000;
            14'h4b14: o_data_a = 16'b1111110111101000;
            14'h4b15: o_data_a = 16'b1110110010100000;
            14'h4b16: o_data_a = 16'b1110001100001000;
            14'h4b17: o_data_a = 16'b0000000000000000;
            14'h4b18: o_data_a = 16'b1111110010101000;
            14'h4b19: o_data_a = 16'b1111110000010000;
            14'h4b1a: o_data_a = 16'b1110110010100000;
            14'h4b1b: o_data_a = 16'b1111000010001000;
            14'h4b1c: o_data_a = 16'b0000000000000001;
            14'h4b1d: o_data_a = 16'b1111110111100000;
            14'h4b1e: o_data_a = 16'b1111110000010000;
            14'h4b1f: o_data_a = 16'b0000000000000000;
            14'h4b20: o_data_a = 16'b1111110111101000;
            14'h4b21: o_data_a = 16'b1110110010100000;
            14'h4b22: o_data_a = 16'b1110001100001000;
            14'h4b23: o_data_a = 16'b0000000000000001;
            14'h4b24: o_data_a = 16'b1111110111100000;
            14'h4b25: o_data_a = 16'b1110110111100000;
            14'h4b26: o_data_a = 16'b1111110000010000;
            14'h4b27: o_data_a = 16'b0000000000000000;
            14'h4b28: o_data_a = 16'b1111110111101000;
            14'h4b29: o_data_a = 16'b1110110010100000;
            14'h4b2a: o_data_a = 16'b1110001100001000;
            14'h4b2b: o_data_a = 16'b0000000000000000;
            14'h4b2c: o_data_a = 16'b1111110010101000;
            14'h4b2d: o_data_a = 16'b1111110000010000;
            14'h4b2e: o_data_a = 16'b1110110010100000;
            14'h4b2f: o_data_a = 16'b1111000010001000;
            14'h4b30: o_data_a = 16'b0000000000000000;
            14'h4b31: o_data_a = 16'b1111110010101000;
            14'h4b32: o_data_a = 16'b1111110000010000;
            14'h4b33: o_data_a = 16'b0000000000000100;
            14'h4b34: o_data_a = 16'b1110001100001000;
            14'h4b35: o_data_a = 16'b0000000000000100;
            14'h4b36: o_data_a = 16'b1111110000100000;
            14'h4b37: o_data_a = 16'b1111110000010000;
            14'h4b38: o_data_a = 16'b0000000000000000;
            14'h4b39: o_data_a = 16'b1111110111101000;
            14'h4b3a: o_data_a = 16'b1110110010100000;
            14'h4b3b: o_data_a = 16'b1110001100001000;
            14'h4b3c: o_data_a = 16'b0000000000000001;
            14'h4b3d: o_data_a = 16'b1111110000010000;
            14'h4b3e: o_data_a = 16'b0000000000000011;
            14'h4b3f: o_data_a = 16'b1110000010100000;
            14'h4b40: o_data_a = 16'b1111110000010000;
            14'h4b41: o_data_a = 16'b0000000000000000;
            14'h4b42: o_data_a = 16'b1111110111101000;
            14'h4b43: o_data_a = 16'b1110110010100000;
            14'h4b44: o_data_a = 16'b1110001100001000;
            14'h4b45: o_data_a = 16'b0000000000000000;
            14'h4b46: o_data_a = 16'b1111110010101000;
            14'h4b47: o_data_a = 16'b1111110000010000;
            14'h4b48: o_data_a = 16'b1110110010100000;
            14'h4b49: o_data_a = 16'b1111010101001000;
            14'h4b4a: o_data_a = 16'b0000000000000000;
            14'h4b4b: o_data_a = 16'b1111110010101000;
            14'h4b4c: o_data_a = 16'b1111110000010000;
            14'h4b4d: o_data_a = 16'b0000000000000101;
            14'h4b4e: o_data_a = 16'b1110001100001000;
            14'h4b4f: o_data_a = 16'b0000000000000000;
            14'h4b50: o_data_a = 16'b1111110010101000;
            14'h4b51: o_data_a = 16'b1111110000010000;
            14'h4b52: o_data_a = 16'b0000000000000100;
            14'h4b53: o_data_a = 16'b1110001100001000;
            14'h4b54: o_data_a = 16'b0000000000000101;
            14'h4b55: o_data_a = 16'b1111110000010000;
            14'h4b56: o_data_a = 16'b0000000000000000;
            14'h4b57: o_data_a = 16'b1111110111101000;
            14'h4b58: o_data_a = 16'b1110110010100000;
            14'h4b59: o_data_a = 16'b1110001100001000;
            14'h4b5a: o_data_a = 16'b0000000000000000;
            14'h4b5b: o_data_a = 16'b1111110010101000;
            14'h4b5c: o_data_a = 16'b1111110000010000;
            14'h4b5d: o_data_a = 16'b0000000000000100;
            14'h4b5e: o_data_a = 16'b1111110000100000;
            14'h4b5f: o_data_a = 16'b1110001100001000;
            14'h4b60: o_data_a = 16'b0000000000000001;
            14'h4b61: o_data_a = 16'b1111110000100000;
            14'h4b62: o_data_a = 16'b1111110000010000;
            14'h4b63: o_data_a = 16'b0000000000000000;
            14'h4b64: o_data_a = 16'b1111110111101000;
            14'h4b65: o_data_a = 16'b1110110010100000;
            14'h4b66: o_data_a = 16'b1110001100001000;
            14'h4b67: o_data_a = 16'b0000000000100000;
            14'h4b68: o_data_a = 16'b1110110000010000;
            14'h4b69: o_data_a = 16'b0000000000000000;
            14'h4b6a: o_data_a = 16'b1111110111101000;
            14'h4b6b: o_data_a = 16'b1110110010100000;
            14'h4b6c: o_data_a = 16'b1110001100001000;
            14'h4b6d: o_data_a = 16'b0000000000000000;
            14'h4b6e: o_data_a = 16'b1111110010101000;
            14'h4b6f: o_data_a = 16'b1111110000010000;
            14'h4b70: o_data_a = 16'b1110110010100000;
            14'h4b71: o_data_a = 16'b1111000010001000;
            14'h4b72: o_data_a = 16'b0000000000000000;
            14'h4b73: o_data_a = 16'b1111110010101000;
            14'h4b74: o_data_a = 16'b1111110000010000;
            14'h4b75: o_data_a = 16'b0000000000000001;
            14'h4b76: o_data_a = 16'b1111110000100000;
            14'h4b77: o_data_a = 16'b1110001100001000;
            14'h4b78: o_data_a = 16'b0000000000000001;
            14'h4b79: o_data_a = 16'b1111110111100000;
            14'h4b7a: o_data_a = 16'b1111110000010000;
            14'h4b7b: o_data_a = 16'b0000000000000000;
            14'h4b7c: o_data_a = 16'b1111110111101000;
            14'h4b7d: o_data_a = 16'b1110110010100000;
            14'h4b7e: o_data_a = 16'b1110001100001000;
            14'h4b7f: o_data_a = 16'b0000000000000000;
            14'h4b80: o_data_a = 16'b1111110111001000;
            14'h4b81: o_data_a = 16'b1111110010100000;
            14'h4b82: o_data_a = 16'b1110111111001000;
            14'h4b83: o_data_a = 16'b0000000000000000;
            14'h4b84: o_data_a = 16'b1111110010101000;
            14'h4b85: o_data_a = 16'b1111110000010000;
            14'h4b86: o_data_a = 16'b1110110010100000;
            14'h4b87: o_data_a = 16'b1111000010001000;
            14'h4b88: o_data_a = 16'b0000000000000000;
            14'h4b89: o_data_a = 16'b1111110010101000;
            14'h4b8a: o_data_a = 16'b1111110000010000;
            14'h4b8b: o_data_a = 16'b0000000000000001;
            14'h4b8c: o_data_a = 16'b1111110111100000;
            14'h4b8d: o_data_a = 16'b1110001100001000;
            14'h4b8e: o_data_a = 16'b0100101001111100;
            14'h4b8f: o_data_a = 16'b1110101010000111;
            14'h4b90: o_data_a = 16'b0000000000000000;
            14'h4b91: o_data_a = 16'b1111110111001000;
            14'h4b92: o_data_a = 16'b1111110010100000;
            14'h4b93: o_data_a = 16'b1110101010001000;
            14'h4b94: o_data_a = 16'b0000000000110110;
            14'h4b95: o_data_a = 16'b1110101010000111;
            14'h4b96: o_data_a = 16'b0000000000000010;
            14'h4b97: o_data_a = 16'b1111110000100000;
            14'h4b98: o_data_a = 16'b1111110000010000;
            14'h4b99: o_data_a = 16'b0000000000000000;
            14'h4b9a: o_data_a = 16'b1111110111101000;
            14'h4b9b: o_data_a = 16'b1110110010100000;
            14'h4b9c: o_data_a = 16'b1110001100001000;
            14'h4b9d: o_data_a = 16'b0000000000000000;
            14'h4b9e: o_data_a = 16'b1111110111001000;
            14'h4b9f: o_data_a = 16'b1111110010100000;
            14'h4ba0: o_data_a = 16'b1110101010001000;
            14'h4ba1: o_data_a = 16'b0100101110100101;
            14'h4ba2: o_data_a = 16'b1110110000010000;
            14'h4ba3: o_data_a = 16'b0000000000100110;
            14'h4ba4: o_data_a = 16'b1110101010000111;
            14'h4ba5: o_data_a = 16'b0000000000000010;
            14'h4ba6: o_data_a = 16'b1111110000100000;
            14'h4ba7: o_data_a = 16'b1111110000010000;
            14'h4ba8: o_data_a = 16'b0000000000000000;
            14'h4ba9: o_data_a = 16'b1111110111101000;
            14'h4baa: o_data_a = 16'b1110110010100000;
            14'h4bab: o_data_a = 16'b1110001100001000;
            14'h4bac: o_data_a = 16'b0000000000010110;
            14'h4bad: o_data_a = 16'b1110110000010000;
            14'h4bae: o_data_a = 16'b0000000000000000;
            14'h4baf: o_data_a = 16'b1111110111101000;
            14'h4bb0: o_data_a = 16'b1110110010100000;
            14'h4bb1: o_data_a = 16'b1110001100001000;
            14'h4bb2: o_data_a = 16'b0100101110110110;
            14'h4bb3: o_data_a = 16'b1110110000010000;
            14'h4bb4: o_data_a = 16'b0000000000010110;
            14'h4bb5: o_data_a = 16'b1110101010000111;
            14'h4bb6: o_data_a = 16'b0000000000000000;
            14'h4bb7: o_data_a = 16'b1111110010101000;
            14'h4bb8: o_data_a = 16'b1111110000010000;
            14'h4bb9: o_data_a = 16'b1110110010100000;
            14'h4bba: o_data_a = 16'b1111010101001000;
            14'h4bbb: o_data_a = 16'b0000000000000010;
            14'h4bbc: o_data_a = 16'b1111110111100000;
            14'h4bbd: o_data_a = 16'b1111110000010000;
            14'h4bbe: o_data_a = 16'b0000000000000000;
            14'h4bbf: o_data_a = 16'b1111110111101000;
            14'h4bc0: o_data_a = 16'b1110110010100000;
            14'h4bc1: o_data_a = 16'b1110001100001000;
            14'h4bc2: o_data_a = 16'b0000000000000000;
            14'h4bc3: o_data_a = 16'b1111110111001000;
            14'h4bc4: o_data_a = 16'b1111110010100000;
            14'h4bc5: o_data_a = 16'b1110101010001000;
            14'h4bc6: o_data_a = 16'b0100101111001010;
            14'h4bc7: o_data_a = 16'b1110110000010000;
            14'h4bc8: o_data_a = 16'b0000000000100110;
            14'h4bc9: o_data_a = 16'b1110101010000111;
            14'h4bca: o_data_a = 16'b0000000000000000;
            14'h4bcb: o_data_a = 16'b1111110010101000;
            14'h4bcc: o_data_a = 16'b1111110000010000;
            14'h4bcd: o_data_a = 16'b1110110010100000;
            14'h4bce: o_data_a = 16'b1111010101001000;
            14'h4bcf: o_data_a = 16'b0000000000000010;
            14'h4bd0: o_data_a = 16'b1111110111100000;
            14'h4bd1: o_data_a = 16'b1111110000010000;
            14'h4bd2: o_data_a = 16'b0000000000000000;
            14'h4bd3: o_data_a = 16'b1111110111101000;
            14'h4bd4: o_data_a = 16'b1110110010100000;
            14'h4bd5: o_data_a = 16'b1110001100001000;
            14'h4bd6: o_data_a = 16'b0000000000111111;
            14'h4bd7: o_data_a = 16'b1110110000010000;
            14'h4bd8: o_data_a = 16'b0000000000000000;
            14'h4bd9: o_data_a = 16'b1111110111101000;
            14'h4bda: o_data_a = 16'b1110110010100000;
            14'h4bdb: o_data_a = 16'b1110001100001000;
            14'h4bdc: o_data_a = 16'b0100101111100000;
            14'h4bdd: o_data_a = 16'b1110110000010000;
            14'h4bde: o_data_a = 16'b0000000000010110;
            14'h4bdf: o_data_a = 16'b1110101010000111;
            14'h4be0: o_data_a = 16'b0000000000000000;
            14'h4be1: o_data_a = 16'b1111110010101000;
            14'h4be2: o_data_a = 16'b1111110000010000;
            14'h4be3: o_data_a = 16'b1110110010100000;
            14'h4be4: o_data_a = 16'b1111010101001000;
            14'h4be5: o_data_a = 16'b0000000000000000;
            14'h4be6: o_data_a = 16'b1111110010101000;
            14'h4be7: o_data_a = 16'b1111110000010000;
            14'h4be8: o_data_a = 16'b0100101111101100;
            14'h4be9: o_data_a = 16'b1110001100000101;
            14'h4bea: o_data_a = 16'b0100110000000011;
            14'h4beb: o_data_a = 16'b1110101010000111;
            14'h4bec: o_data_a = 16'b0000000000010100;
            14'h4bed: o_data_a = 16'b1110110000010000;
            14'h4bee: o_data_a = 16'b0000000000000000;
            14'h4bef: o_data_a = 16'b1111110111101000;
            14'h4bf0: o_data_a = 16'b1110110010100000;
            14'h4bf1: o_data_a = 16'b1110001100001000;
            14'h4bf2: o_data_a = 16'b0000000000000001;
            14'h4bf3: o_data_a = 16'b1110110000010000;
            14'h4bf4: o_data_a = 16'b0000000000001101;
            14'h4bf5: o_data_a = 16'b1110001100001000;
            14'h4bf6: o_data_a = 16'b0110101011011001;
            14'h4bf7: o_data_a = 16'b1110110000010000;
            14'h4bf8: o_data_a = 16'b0000000000001110;
            14'h4bf9: o_data_a = 16'b1110001100001000;
            14'h4bfa: o_data_a = 16'b0100101111111110;
            14'h4bfb: o_data_a = 16'b1110110000010000;
            14'h4bfc: o_data_a = 16'b0000000001011111;
            14'h4bfd: o_data_a = 16'b1110101010000111;
            14'h4bfe: o_data_a = 16'b0000000000000000;
            14'h4bff: o_data_a = 16'b1111110010101000;
            14'h4c00: o_data_a = 16'b1111110000010000;
            14'h4c01: o_data_a = 16'b0000000000000101;
            14'h4c02: o_data_a = 16'b1110001100001000;
            14'h4c03: o_data_a = 16'b0000000000000010;
            14'h4c04: o_data_a = 16'b1111110111100000;
            14'h4c05: o_data_a = 16'b1111110000010000;
            14'h4c06: o_data_a = 16'b0000000000000000;
            14'h4c07: o_data_a = 16'b1111110111101000;
            14'h4c08: o_data_a = 16'b1110110010100000;
            14'h4c09: o_data_a = 16'b1110001100001000;
            14'h4c0a: o_data_a = 16'b0000000000000010;
            14'h4c0b: o_data_a = 16'b1110110000010000;
            14'h4c0c: o_data_a = 16'b0000000000000000;
            14'h4c0d: o_data_a = 16'b1111110111101000;
            14'h4c0e: o_data_a = 16'b1110110010100000;
            14'h4c0f: o_data_a = 16'b1110001100001000;
            14'h4c10: o_data_a = 16'b0000000000000010;
            14'h4c11: o_data_a = 16'b1110110000010000;
            14'h4c12: o_data_a = 16'b0000000000001101;
            14'h4c13: o_data_a = 16'b1110001100001000;
            14'h4c14: o_data_a = 16'b0001110001110111;
            14'h4c15: o_data_a = 16'b1110110000010000;
            14'h4c16: o_data_a = 16'b0000000000001110;
            14'h4c17: o_data_a = 16'b1110001100001000;
            14'h4c18: o_data_a = 16'b0100110000011100;
            14'h4c19: o_data_a = 16'b1110110000010000;
            14'h4c1a: o_data_a = 16'b0000000001011111;
            14'h4c1b: o_data_a = 16'b1110101010000111;
            14'h4c1c: o_data_a = 16'b0000000000000000;
            14'h4c1d: o_data_a = 16'b1111110010101000;
            14'h4c1e: o_data_a = 16'b1111110000010000;
            14'h4c1f: o_data_a = 16'b0000000000010111;
            14'h4c20: o_data_a = 16'b1110001100001000;
            14'h4c21: o_data_a = 16'b0000000000100000;
            14'h4c22: o_data_a = 16'b1110110000010000;
            14'h4c23: o_data_a = 16'b0000000000000000;
            14'h4c24: o_data_a = 16'b1111110111101000;
            14'h4c25: o_data_a = 16'b1110110010100000;
            14'h4c26: o_data_a = 16'b1110001100001000;
            14'h4c27: o_data_a = 16'b0000000000000010;
            14'h4c28: o_data_a = 16'b1111110000100000;
            14'h4c29: o_data_a = 16'b1111110000010000;
            14'h4c2a: o_data_a = 16'b0000000000000000;
            14'h4c2b: o_data_a = 16'b1111110111101000;
            14'h4c2c: o_data_a = 16'b1110110010100000;
            14'h4c2d: o_data_a = 16'b1110001100001000;
            14'h4c2e: o_data_a = 16'b0000000101100000;
            14'h4c2f: o_data_a = 16'b1110110000010000;
            14'h4c30: o_data_a = 16'b0000000000000000;
            14'h4c31: o_data_a = 16'b1111110111101000;
            14'h4c32: o_data_a = 16'b1110110010100000;
            14'h4c33: o_data_a = 16'b1110001100001000;
            14'h4c34: o_data_a = 16'b0000000000000010;
            14'h4c35: o_data_a = 16'b1110110000010000;
            14'h4c36: o_data_a = 16'b0000000000001101;
            14'h4c37: o_data_a = 16'b1110001100001000;
            14'h4c38: o_data_a = 16'b0001101010100110;
            14'h4c39: o_data_a = 16'b1110110000010000;
            14'h4c3a: o_data_a = 16'b0000000000001110;
            14'h4c3b: o_data_a = 16'b1110001100001000;
            14'h4c3c: o_data_a = 16'b0100110001000000;
            14'h4c3d: o_data_a = 16'b1110110000010000;
            14'h4c3e: o_data_a = 16'b0000000001011111;
            14'h4c3f: o_data_a = 16'b1110101010000111;
            14'h4c40: o_data_a = 16'b0000000000000000;
            14'h4c41: o_data_a = 16'b1111110010101000;
            14'h4c42: o_data_a = 16'b1111110000010000;
            14'h4c43: o_data_a = 16'b1110110010100000;
            14'h4c44: o_data_a = 16'b1111000010001000;
            14'h4c45: o_data_a = 16'b0000000000010111;
            14'h4c46: o_data_a = 16'b1111110000010000;
            14'h4c47: o_data_a = 16'b0000000000000000;
            14'h4c48: o_data_a = 16'b1111110111101000;
            14'h4c49: o_data_a = 16'b1110110010100000;
            14'h4c4a: o_data_a = 16'b1110001100001000;
            14'h4c4b: o_data_a = 16'b0000000000000000;
            14'h4c4c: o_data_a = 16'b1111110010101000;
            14'h4c4d: o_data_a = 16'b1111110000010000;
            14'h4c4e: o_data_a = 16'b1110110010100000;
            14'h4c4f: o_data_a = 16'b1111000010001000;
            14'h4c50: o_data_a = 16'b0000000000000000;
            14'h4c51: o_data_a = 16'b1111110010101000;
            14'h4c52: o_data_a = 16'b1111110000010000;
            14'h4c53: o_data_a = 16'b0000000000010110;
            14'h4c54: o_data_a = 16'b1110001100001000;
            14'h4c55: o_data_a = 16'b0000000000000010;
            14'h4c56: o_data_a = 16'b1111110111100000;
            14'h4c57: o_data_a = 16'b1111110000010000;
            14'h4c58: o_data_a = 16'b0000000000000000;
            14'h4c59: o_data_a = 16'b1111110111101000;
            14'h4c5a: o_data_a = 16'b1110110010100000;
            14'h4c5b: o_data_a = 16'b1110001100001000;
            14'h4c5c: o_data_a = 16'b0000000000010111;
            14'h4c5d: o_data_a = 16'b1111110000010000;
            14'h4c5e: o_data_a = 16'b0000000000000000;
            14'h4c5f: o_data_a = 16'b1111110111101000;
            14'h4c60: o_data_a = 16'b1110110010100000;
            14'h4c61: o_data_a = 16'b1110001100001000;
            14'h4c62: o_data_a = 16'b0000000000000010;
            14'h4c63: o_data_a = 16'b1110110000010000;
            14'h4c64: o_data_a = 16'b0000000000000000;
            14'h4c65: o_data_a = 16'b1111110111101000;
            14'h4c66: o_data_a = 16'b1110110010100000;
            14'h4c67: o_data_a = 16'b1110001100001000;
            14'h4c68: o_data_a = 16'b0000000000000010;
            14'h4c69: o_data_a = 16'b1110110000010000;
            14'h4c6a: o_data_a = 16'b0000000000001101;
            14'h4c6b: o_data_a = 16'b1110001100001000;
            14'h4c6c: o_data_a = 16'b0001101010100110;
            14'h4c6d: o_data_a = 16'b1110110000010000;
            14'h4c6e: o_data_a = 16'b0000000000001110;
            14'h4c6f: o_data_a = 16'b1110001100001000;
            14'h4c70: o_data_a = 16'b0100110001110100;
            14'h4c71: o_data_a = 16'b1110110000010000;
            14'h4c72: o_data_a = 16'b0000000001011111;
            14'h4c73: o_data_a = 16'b1110101010000111;
            14'h4c74: o_data_a = 16'b0100110001111000;
            14'h4c75: o_data_a = 16'b1110110000010000;
            14'h4c76: o_data_a = 16'b0000000000000110;
            14'h4c77: o_data_a = 16'b1110101010000111;
            14'h4c78: o_data_a = 16'b0000000000000000;
            14'h4c79: o_data_a = 16'b1111110010101000;
            14'h4c7a: o_data_a = 16'b1111110000010000;
            14'h4c7b: o_data_a = 16'b0000000000010101;
            14'h4c7c: o_data_a = 16'b1110001100001000;
            14'h4c7d: o_data_a = 16'b0000000000100000;
            14'h4c7e: o_data_a = 16'b1110110000010000;
            14'h4c7f: o_data_a = 16'b0000000000000000;
            14'h4c80: o_data_a = 16'b1111110111101000;
            14'h4c81: o_data_a = 16'b1110110010100000;
            14'h4c82: o_data_a = 16'b1110001100001000;
            14'h4c83: o_data_a = 16'b0000000000000001;
            14'h4c84: o_data_a = 16'b1110110000010000;
            14'h4c85: o_data_a = 16'b0000000000001101;
            14'h4c86: o_data_a = 16'b1110001100001000;
            14'h4c87: o_data_a = 16'b0100101001001101;
            14'h4c88: o_data_a = 16'b1110110000010000;
            14'h4c89: o_data_a = 16'b0000000000001110;
            14'h4c8a: o_data_a = 16'b1110001100001000;
            14'h4c8b: o_data_a = 16'b0100110010001111;
            14'h4c8c: o_data_a = 16'b1110110000010000;
            14'h4c8d: o_data_a = 16'b0000000001011111;
            14'h4c8e: o_data_a = 16'b1110101010000111;
            14'h4c8f: o_data_a = 16'b0000000000000000;
            14'h4c90: o_data_a = 16'b1111110010101000;
            14'h4c91: o_data_a = 16'b1111110000010000;
            14'h4c92: o_data_a = 16'b0000000000000101;
            14'h4c93: o_data_a = 16'b1110001100001000;
            14'h4c94: o_data_a = 16'b0000000000000000;
            14'h4c95: o_data_a = 16'b1111110111001000;
            14'h4c96: o_data_a = 16'b1111110010100000;
            14'h4c97: o_data_a = 16'b1110101010001000;
            14'h4c98: o_data_a = 16'b0000000000110110;
            14'h4c99: o_data_a = 16'b1110101010000111;
            14'h4c9a: o_data_a = 16'b0000000000000010;
            14'h4c9b: o_data_a = 16'b1111110000100000;
            14'h4c9c: o_data_a = 16'b1111110000010000;
            14'h4c9d: o_data_a = 16'b0000000000000000;
            14'h4c9e: o_data_a = 16'b1111110111101000;
            14'h4c9f: o_data_a = 16'b1110110010100000;
            14'h4ca0: o_data_a = 16'b1110001100001000;
            14'h4ca1: o_data_a = 16'b0000000000000000;
            14'h4ca2: o_data_a = 16'b1110110000010000;
            14'h4ca3: o_data_a = 16'b0000000000001101;
            14'h4ca4: o_data_a = 16'b1110001100001000;
            14'h4ca5: o_data_a = 16'b0110100110011010;
            14'h4ca6: o_data_a = 16'b1110110000010000;
            14'h4ca7: o_data_a = 16'b0000000000001110;
            14'h4ca8: o_data_a = 16'b1110001100001000;
            14'h4ca9: o_data_a = 16'b0100110010101101;
            14'h4caa: o_data_a = 16'b1110110000010000;
            14'h4cab: o_data_a = 16'b0000000001011111;
            14'h4cac: o_data_a = 16'b1110101010000111;
            14'h4cad: o_data_a = 16'b0100110010110001;
            14'h4cae: o_data_a = 16'b1110110000010000;
            14'h4caf: o_data_a = 16'b0000000000000110;
            14'h4cb0: o_data_a = 16'b1110101010000111;
            14'h4cb1: o_data_a = 16'b0000000000000000;
            14'h4cb2: o_data_a = 16'b1111110010101000;
            14'h4cb3: o_data_a = 16'b1111110000010000;
            14'h4cb4: o_data_a = 16'b0100110010111000;
            14'h4cb5: o_data_a = 16'b1110001100000101;
            14'h4cb6: o_data_a = 16'b0100110011001011;
            14'h4cb7: o_data_a = 16'b1110101010000111;
            14'h4cb8: o_data_a = 16'b0000000000000000;
            14'h4cb9: o_data_a = 16'b1110110000010000;
            14'h4cba: o_data_a = 16'b0000000000001101;
            14'h4cbb: o_data_a = 16'b1110001100001000;
            14'h4cbc: o_data_a = 16'b0100111001001000;
            14'h4cbd: o_data_a = 16'b1110110000010000;
            14'h4cbe: o_data_a = 16'b0000000000001110;
            14'h4cbf: o_data_a = 16'b1110001100001000;
            14'h4cc0: o_data_a = 16'b0100110011000100;
            14'h4cc1: o_data_a = 16'b1110110000010000;
            14'h4cc2: o_data_a = 16'b0000000001011111;
            14'h4cc3: o_data_a = 16'b1110101010000111;
            14'h4cc4: o_data_a = 16'b0000000000000000;
            14'h4cc5: o_data_a = 16'b1111110010101000;
            14'h4cc6: o_data_a = 16'b1111110000010000;
            14'h4cc7: o_data_a = 16'b0000000000000101;
            14'h4cc8: o_data_a = 16'b1110001100001000;
            14'h4cc9: o_data_a = 16'b0100110110000100;
            14'h4cca: o_data_a = 16'b1110101010000111;
            14'h4ccb: o_data_a = 16'b0000000000000010;
            14'h4ccc: o_data_a = 16'b1111110000100000;
            14'h4ccd: o_data_a = 16'b1111110000010000;
            14'h4cce: o_data_a = 16'b0000000000000000;
            14'h4ccf: o_data_a = 16'b1111110111101000;
            14'h4cd0: o_data_a = 16'b1110110010100000;
            14'h4cd1: o_data_a = 16'b1110001100001000;
            14'h4cd2: o_data_a = 16'b0000000000000000;
            14'h4cd3: o_data_a = 16'b1110110000010000;
            14'h4cd4: o_data_a = 16'b0000000000001101;
            14'h4cd5: o_data_a = 16'b1110001100001000;
            14'h4cd6: o_data_a = 16'b0110100110100010;
            14'h4cd7: o_data_a = 16'b1110110000010000;
            14'h4cd8: o_data_a = 16'b0000000000001110;
            14'h4cd9: o_data_a = 16'b1110001100001000;
            14'h4cda: o_data_a = 16'b0100110011011110;
            14'h4cdb: o_data_a = 16'b1110110000010000;
            14'h4cdc: o_data_a = 16'b0000000001011111;
            14'h4cdd: o_data_a = 16'b1110101010000111;
            14'h4cde: o_data_a = 16'b0100110011100010;
            14'h4cdf: o_data_a = 16'b1110110000010000;
            14'h4ce0: o_data_a = 16'b0000000000000110;
            14'h4ce1: o_data_a = 16'b1110101010000111;
            14'h4ce2: o_data_a = 16'b0000000000000000;
            14'h4ce3: o_data_a = 16'b1111110010101000;
            14'h4ce4: o_data_a = 16'b1111110000010000;
            14'h4ce5: o_data_a = 16'b0100110011101001;
            14'h4ce6: o_data_a = 16'b1110001100000101;
            14'h4ce7: o_data_a = 16'b0100110011111100;
            14'h4ce8: o_data_a = 16'b1110101010000111;
            14'h4ce9: o_data_a = 16'b0000000000000000;
            14'h4cea: o_data_a = 16'b1110110000010000;
            14'h4ceb: o_data_a = 16'b0000000000001101;
            14'h4cec: o_data_a = 16'b1110001100001000;
            14'h4ced: o_data_a = 16'b0100111010100110;
            14'h4cee: o_data_a = 16'b1110110000010000;
            14'h4cef: o_data_a = 16'b0000000000001110;
            14'h4cf0: o_data_a = 16'b1110001100001000;
            14'h4cf1: o_data_a = 16'b0100110011110101;
            14'h4cf2: o_data_a = 16'b1110110000010000;
            14'h4cf3: o_data_a = 16'b0000000001011111;
            14'h4cf4: o_data_a = 16'b1110101010000111;
            14'h4cf5: o_data_a = 16'b0000000000000000;
            14'h4cf6: o_data_a = 16'b1111110010101000;
            14'h4cf7: o_data_a = 16'b1111110000010000;
            14'h4cf8: o_data_a = 16'b0000000000000101;
            14'h4cf9: o_data_a = 16'b1110001100001000;
            14'h4cfa: o_data_a = 16'b0100110110000100;
            14'h4cfb: o_data_a = 16'b1110101010000111;
            14'h4cfc: o_data_a = 16'b0000000000000010;
            14'h4cfd: o_data_a = 16'b1111110000100000;
            14'h4cfe: o_data_a = 16'b1111110000010000;
            14'h4cff: o_data_a = 16'b0000000000000000;
            14'h4d00: o_data_a = 16'b1111110111101000;
            14'h4d01: o_data_a = 16'b1110110010100000;
            14'h4d02: o_data_a = 16'b1110001100001000;
            14'h4d03: o_data_a = 16'b0000000000000001;
            14'h4d04: o_data_a = 16'b1110110000010000;
            14'h4d05: o_data_a = 16'b0000000000001101;
            14'h4d06: o_data_a = 16'b1110001100001000;
            14'h4d07: o_data_a = 16'b0100101001001101;
            14'h4d08: o_data_a = 16'b1110110000010000;
            14'h4d09: o_data_a = 16'b0000000000001110;
            14'h4d0a: o_data_a = 16'b1110001100001000;
            14'h4d0b: o_data_a = 16'b0100110100001111;
            14'h4d0c: o_data_a = 16'b1110110000010000;
            14'h4d0d: o_data_a = 16'b0000000001011111;
            14'h4d0e: o_data_a = 16'b1110101010000111;
            14'h4d0f: o_data_a = 16'b0000000000000000;
            14'h4d10: o_data_a = 16'b1111110010101000;
            14'h4d11: o_data_a = 16'b1111110000010000;
            14'h4d12: o_data_a = 16'b0000000000000101;
            14'h4d13: o_data_a = 16'b1110001100001000;
            14'h4d14: o_data_a = 16'b0000000000010101;
            14'h4d15: o_data_a = 16'b1111110000010000;
            14'h4d16: o_data_a = 16'b0000000000000000;
            14'h4d17: o_data_a = 16'b1111110111101000;
            14'h4d18: o_data_a = 16'b1110110010100000;
            14'h4d19: o_data_a = 16'b1110001100001000;
            14'h4d1a: o_data_a = 16'b0000000000000000;
            14'h4d1b: o_data_a = 16'b1111110010100000;
            14'h4d1c: o_data_a = 16'b1111110001001000;
            14'h4d1d: o_data_a = 16'b0000000000000000;
            14'h4d1e: o_data_a = 16'b1111110010101000;
            14'h4d1f: o_data_a = 16'b1111110000010000;
            14'h4d20: o_data_a = 16'b0100110100100100;
            14'h4d21: o_data_a = 16'b1110001100000101;
            14'h4d22: o_data_a = 16'b0100110101001100;
            14'h4d23: o_data_a = 16'b1110101010000111;
            14'h4d24: o_data_a = 16'b0000000000010111;
            14'h4d25: o_data_a = 16'b1111110000010000;
            14'h4d26: o_data_a = 16'b0000000000000000;
            14'h4d27: o_data_a = 16'b1111110111101000;
            14'h4d28: o_data_a = 16'b1110110010100000;
            14'h4d29: o_data_a = 16'b1110001100001000;
            14'h4d2a: o_data_a = 16'b0000000000000000;
            14'h4d2b: o_data_a = 16'b1111110111001000;
            14'h4d2c: o_data_a = 16'b1111110010100000;
            14'h4d2d: o_data_a = 16'b1110111111001000;
            14'h4d2e: o_data_a = 16'b0000000000000000;
            14'h4d2f: o_data_a = 16'b1111110010101000;
            14'h4d30: o_data_a = 16'b1111110000010000;
            14'h4d31: o_data_a = 16'b1110110010100000;
            14'h4d32: o_data_a = 16'b1111000010001000;
            14'h4d33: o_data_a = 16'b0000000000000000;
            14'h4d34: o_data_a = 16'b1111110010101000;
            14'h4d35: o_data_a = 16'b1111110000010000;
            14'h4d36: o_data_a = 16'b0000000000010111;
            14'h4d37: o_data_a = 16'b1110001100001000;
            14'h4d38: o_data_a = 16'b0000000000010110;
            14'h4d39: o_data_a = 16'b1111110000010000;
            14'h4d3a: o_data_a = 16'b0000000000000000;
            14'h4d3b: o_data_a = 16'b1111110111101000;
            14'h4d3c: o_data_a = 16'b1110110010100000;
            14'h4d3d: o_data_a = 16'b1110001100001000;
            14'h4d3e: o_data_a = 16'b0000000000000000;
            14'h4d3f: o_data_a = 16'b1111110111001000;
            14'h4d40: o_data_a = 16'b1111110010100000;
            14'h4d41: o_data_a = 16'b1110111111001000;
            14'h4d42: o_data_a = 16'b0000000000000000;
            14'h4d43: o_data_a = 16'b1111110010101000;
            14'h4d44: o_data_a = 16'b1111110000010000;
            14'h4d45: o_data_a = 16'b1110110010100000;
            14'h4d46: o_data_a = 16'b1111000010001000;
            14'h4d47: o_data_a = 16'b0000000000000000;
            14'h4d48: o_data_a = 16'b1111110010101000;
            14'h4d49: o_data_a = 16'b1111110000010000;
            14'h4d4a: o_data_a = 16'b0000000000010110;
            14'h4d4b: o_data_a = 16'b1110001100001000;
            14'h4d4c: o_data_a = 16'b0000000000010111;
            14'h4d4d: o_data_a = 16'b1111110000010000;
            14'h4d4e: o_data_a = 16'b0000000000000000;
            14'h4d4f: o_data_a = 16'b1111110111101000;
            14'h4d50: o_data_a = 16'b1110110010100000;
            14'h4d51: o_data_a = 16'b1110001100001000;
            14'h4d52: o_data_a = 16'b0000000000100000;
            14'h4d53: o_data_a = 16'b1110110000010000;
            14'h4d54: o_data_a = 16'b0000000000000000;
            14'h4d55: o_data_a = 16'b1111110111101000;
            14'h4d56: o_data_a = 16'b1110110010100000;
            14'h4d57: o_data_a = 16'b1110001100001000;
            14'h4d58: o_data_a = 16'b0100110101011100;
            14'h4d59: o_data_a = 16'b1110110000010000;
            14'h4d5a: o_data_a = 16'b0000000000000110;
            14'h4d5b: o_data_a = 16'b1110101010000111;
            14'h4d5c: o_data_a = 16'b0000000000000000;
            14'h4d5d: o_data_a = 16'b1111110010101000;
            14'h4d5e: o_data_a = 16'b1111110000010000;
            14'h4d5f: o_data_a = 16'b0100110101100011;
            14'h4d60: o_data_a = 16'b1110001100000101;
            14'h4d61: o_data_a = 16'b0100110101110110;
            14'h4d62: o_data_a = 16'b1110101010000111;
            14'h4d63: o_data_a = 16'b0000000000000000;
            14'h4d64: o_data_a = 16'b1110110000010000;
            14'h4d65: o_data_a = 16'b0000000000001101;
            14'h4d66: o_data_a = 16'b1110001100001000;
            14'h4d67: o_data_a = 16'b0100111001001000;
            14'h4d68: o_data_a = 16'b1110110000010000;
            14'h4d69: o_data_a = 16'b0000000000001110;
            14'h4d6a: o_data_a = 16'b1110001100001000;
            14'h4d6b: o_data_a = 16'b0100110101101111;
            14'h4d6c: o_data_a = 16'b1110110000010000;
            14'h4d6d: o_data_a = 16'b0000000001011111;
            14'h4d6e: o_data_a = 16'b1110101010000111;
            14'h4d6f: o_data_a = 16'b0000000000000000;
            14'h4d70: o_data_a = 16'b1111110010101000;
            14'h4d71: o_data_a = 16'b1111110000010000;
            14'h4d72: o_data_a = 16'b0000000000000101;
            14'h4d73: o_data_a = 16'b1110001100001000;
            14'h4d74: o_data_a = 16'b0100110110000100;
            14'h4d75: o_data_a = 16'b1110101010000111;
            14'h4d76: o_data_a = 16'b0000000000010101;
            14'h4d77: o_data_a = 16'b1111110000010000;
            14'h4d78: o_data_a = 16'b0000000000000000;
            14'h4d79: o_data_a = 16'b1111110111101000;
            14'h4d7a: o_data_a = 16'b1110110010100000;
            14'h4d7b: o_data_a = 16'b1110001100001000;
            14'h4d7c: o_data_a = 16'b0000000000000000;
            14'h4d7d: o_data_a = 16'b1111110010100000;
            14'h4d7e: o_data_a = 16'b1111110001001000;
            14'h4d7f: o_data_a = 16'b0000000000000000;
            14'h4d80: o_data_a = 16'b1111110010101000;
            14'h4d81: o_data_a = 16'b1111110000010000;
            14'h4d82: o_data_a = 16'b0000000000010101;
            14'h4d83: o_data_a = 16'b1110001100001000;
            14'h4d84: o_data_a = 16'b0000000000000000;
            14'h4d85: o_data_a = 16'b1111110111001000;
            14'h4d86: o_data_a = 16'b1111110010100000;
            14'h4d87: o_data_a = 16'b1110101010001000;
            14'h4d88: o_data_a = 16'b0000000000110110;
            14'h4d89: o_data_a = 16'b1110101010000111;
            14'h4d8a: o_data_a = 16'b0000000000000000;
            14'h4d8b: o_data_a = 16'b1111110000100000;
            14'h4d8c: o_data_a = 16'b1110101010001000;
            14'h4d8d: o_data_a = 16'b1110110111110000;
            14'h4d8e: o_data_a = 16'b1110101010001000;
            14'h4d8f: o_data_a = 16'b0000000000000000;
            14'h4d90: o_data_a = 16'b1110011111001000;
            14'h4d91: o_data_a = 16'b0000000000000010;
            14'h4d92: o_data_a = 16'b1111110000100000;
            14'h4d93: o_data_a = 16'b1111110000010000;
            14'h4d94: o_data_a = 16'b0000000000000000;
            14'h4d95: o_data_a = 16'b1111110111101000;
            14'h4d96: o_data_a = 16'b1110110010100000;
            14'h4d97: o_data_a = 16'b1110001100001000;
            14'h4d98: o_data_a = 16'b0000000000000001;
            14'h4d99: o_data_a = 16'b1110110000010000;
            14'h4d9a: o_data_a = 16'b0000000000001101;
            14'h4d9b: o_data_a = 16'b1110001100001000;
            14'h4d9c: o_data_a = 16'b0110001011111011;
            14'h4d9d: o_data_a = 16'b1110110000010000;
            14'h4d9e: o_data_a = 16'b0000000000001110;
            14'h4d9f: o_data_a = 16'b1110001100001000;
            14'h4da0: o_data_a = 16'b0100110110100100;
            14'h4da1: o_data_a = 16'b1110110000010000;
            14'h4da2: o_data_a = 16'b0000000001011111;
            14'h4da3: o_data_a = 16'b1110101010000111;
            14'h4da4: o_data_a = 16'b0000000000000000;
            14'h4da5: o_data_a = 16'b1111110010101000;
            14'h4da6: o_data_a = 16'b1111110000010000;
            14'h4da7: o_data_a = 16'b0000000000000001;
            14'h4da8: o_data_a = 16'b1111110111100000;
            14'h4da9: o_data_a = 16'b1110001100001000;
            14'h4daa: o_data_a = 16'b0000000000000001;
            14'h4dab: o_data_a = 16'b1111110000100000;
            14'h4dac: o_data_a = 16'b1111110000010000;
            14'h4dad: o_data_a = 16'b0000000000000000;
            14'h4dae: o_data_a = 16'b1111110111101000;
            14'h4daf: o_data_a = 16'b1110110010100000;
            14'h4db0: o_data_a = 16'b1110001100001000;
            14'h4db1: o_data_a = 16'b0000000000000001;
            14'h4db2: o_data_a = 16'b1111110111100000;
            14'h4db3: o_data_a = 16'b1111110000010000;
            14'h4db4: o_data_a = 16'b0000000000000000;
            14'h4db5: o_data_a = 16'b1111110111101000;
            14'h4db6: o_data_a = 16'b1110110010100000;
            14'h4db7: o_data_a = 16'b1110001100001000;
            14'h4db8: o_data_a = 16'b0100110110111100;
            14'h4db9: o_data_a = 16'b1110110000010000;
            14'h4dba: o_data_a = 16'b0000000000100110;
            14'h4dbb: o_data_a = 16'b1110101010000111;
            14'h4dbc: o_data_a = 16'b0000000000000000;
            14'h4dbd: o_data_a = 16'b1111110010100000;
            14'h4dbe: o_data_a = 16'b1111110001001000;
            14'h4dbf: o_data_a = 16'b0000000000000000;
            14'h4dc0: o_data_a = 16'b1111110010101000;
            14'h4dc1: o_data_a = 16'b1111110000010000;
            14'h4dc2: o_data_a = 16'b0100111000000111;
            14'h4dc3: o_data_a = 16'b1110001100000101;
            14'h4dc4: o_data_a = 16'b0000000000000010;
            14'h4dc5: o_data_a = 16'b1111110000100000;
            14'h4dc6: o_data_a = 16'b1111110000010000;
            14'h4dc7: o_data_a = 16'b0000000000000000;
            14'h4dc8: o_data_a = 16'b1111110111101000;
            14'h4dc9: o_data_a = 16'b1110110010100000;
            14'h4dca: o_data_a = 16'b1110001100001000;
            14'h4dcb: o_data_a = 16'b0000000000000001;
            14'h4dcc: o_data_a = 16'b1111110000100000;
            14'h4dcd: o_data_a = 16'b1111110000010000;
            14'h4dce: o_data_a = 16'b0000000000000000;
            14'h4dcf: o_data_a = 16'b1111110111101000;
            14'h4dd0: o_data_a = 16'b1110110010100000;
            14'h4dd1: o_data_a = 16'b1110001100001000;
            14'h4dd2: o_data_a = 16'b0000000000000010;
            14'h4dd3: o_data_a = 16'b1110110000010000;
            14'h4dd4: o_data_a = 16'b0000000000001101;
            14'h4dd5: o_data_a = 16'b1110001100001000;
            14'h4dd6: o_data_a = 16'b0110001100010001;
            14'h4dd7: o_data_a = 16'b1110110000010000;
            14'h4dd8: o_data_a = 16'b0000000000001110;
            14'h4dd9: o_data_a = 16'b1110001100001000;
            14'h4dda: o_data_a = 16'b0100110111011110;
            14'h4ddb: o_data_a = 16'b1110110000010000;
            14'h4ddc: o_data_a = 16'b0000000001011111;
            14'h4ddd: o_data_a = 16'b1110101010000111;
            14'h4dde: o_data_a = 16'b0000000000000001;
            14'h4ddf: o_data_a = 16'b1110110000010000;
            14'h4de0: o_data_a = 16'b0000000000001101;
            14'h4de1: o_data_a = 16'b1110001100001000;
            14'h4de2: o_data_a = 16'b0100110010011010;
            14'h4de3: o_data_a = 16'b1110110000010000;
            14'h4de4: o_data_a = 16'b0000000000001110;
            14'h4de5: o_data_a = 16'b1110001100001000;
            14'h4de6: o_data_a = 16'b0100110111101010;
            14'h4de7: o_data_a = 16'b1110110000010000;
            14'h4de8: o_data_a = 16'b0000000001011111;
            14'h4de9: o_data_a = 16'b1110101010000111;
            14'h4dea: o_data_a = 16'b0000000000000000;
            14'h4deb: o_data_a = 16'b1111110010101000;
            14'h4dec: o_data_a = 16'b1111110000010000;
            14'h4ded: o_data_a = 16'b0000000000000101;
            14'h4dee: o_data_a = 16'b1110001100001000;
            14'h4def: o_data_a = 16'b0000000000000001;
            14'h4df0: o_data_a = 16'b1111110000100000;
            14'h4df1: o_data_a = 16'b1111110000010000;
            14'h4df2: o_data_a = 16'b0000000000000000;
            14'h4df3: o_data_a = 16'b1111110111101000;
            14'h4df4: o_data_a = 16'b1110110010100000;
            14'h4df5: o_data_a = 16'b1110001100001000;
            14'h4df6: o_data_a = 16'b0000000000000000;
            14'h4df7: o_data_a = 16'b1111110111001000;
            14'h4df8: o_data_a = 16'b1111110010100000;
            14'h4df9: o_data_a = 16'b1110111111001000;
            14'h4dfa: o_data_a = 16'b0000000000000000;
            14'h4dfb: o_data_a = 16'b1111110010101000;
            14'h4dfc: o_data_a = 16'b1111110000010000;
            14'h4dfd: o_data_a = 16'b1110110010100000;
            14'h4dfe: o_data_a = 16'b1111000010001000;
            14'h4dff: o_data_a = 16'b0000000000000000;
            14'h4e00: o_data_a = 16'b1111110010101000;
            14'h4e01: o_data_a = 16'b1111110000010000;
            14'h4e02: o_data_a = 16'b0000000000000001;
            14'h4e03: o_data_a = 16'b1111110000100000;
            14'h4e04: o_data_a = 16'b1110001100001000;
            14'h4e05: o_data_a = 16'b0100110110101010;
            14'h4e06: o_data_a = 16'b1110101010000111;
            14'h4e07: o_data_a = 16'b0000000000000000;
            14'h4e08: o_data_a = 16'b1111110111001000;
            14'h4e09: o_data_a = 16'b1111110010100000;
            14'h4e0a: o_data_a = 16'b1110101010001000;
            14'h4e0b: o_data_a = 16'b0000000000110110;
            14'h4e0c: o_data_a = 16'b1110101010000111;
            14'h4e0d: o_data_a = 16'b0000000000011000;
            14'h4e0e: o_data_a = 16'b1111110000010000;
            14'h4e0f: o_data_a = 16'b0000000000000000;
            14'h4e10: o_data_a = 16'b1111110111101000;
            14'h4e11: o_data_a = 16'b1110110010100000;
            14'h4e12: o_data_a = 16'b1110001100001000;
            14'h4e13: o_data_a = 16'b0000000000000010;
            14'h4e14: o_data_a = 16'b1111110000100000;
            14'h4e15: o_data_a = 16'b1111110000010000;
            14'h4e16: o_data_a = 16'b0000000000000000;
            14'h4e17: o_data_a = 16'b1111110111101000;
            14'h4e18: o_data_a = 16'b1110110010100000;
            14'h4e19: o_data_a = 16'b1110001100001000;
            14'h4e1a: o_data_a = 16'b0000000000000010;
            14'h4e1b: o_data_a = 16'b1110110000010000;
            14'h4e1c: o_data_a = 16'b0000000000001101;
            14'h4e1d: o_data_a = 16'b1110001100001000;
            14'h4e1e: o_data_a = 16'b0110011010110011;
            14'h4e1f: o_data_a = 16'b1110110000010000;
            14'h4e20: o_data_a = 16'b0000000000001110;
            14'h4e21: o_data_a = 16'b1110001100001000;
            14'h4e22: o_data_a = 16'b0100111000100110;
            14'h4e23: o_data_a = 16'b1110110000010000;
            14'h4e24: o_data_a = 16'b0000000001011111;
            14'h4e25: o_data_a = 16'b1110101010000111;
            14'h4e26: o_data_a = 16'b0000000000000000;
            14'h4e27: o_data_a = 16'b1111110010101000;
            14'h4e28: o_data_a = 16'b1111110000010000;
            14'h4e29: o_data_a = 16'b0000000000000101;
            14'h4e2a: o_data_a = 16'b1110001100001000;
            14'h4e2b: o_data_a = 16'b0000000000011000;
            14'h4e2c: o_data_a = 16'b1111110000010000;
            14'h4e2d: o_data_a = 16'b0000000000000000;
            14'h4e2e: o_data_a = 16'b1111110111101000;
            14'h4e2f: o_data_a = 16'b1110110010100000;
            14'h4e30: o_data_a = 16'b1110001100001000;
            14'h4e31: o_data_a = 16'b0000000000000001;
            14'h4e32: o_data_a = 16'b1110110000010000;
            14'h4e33: o_data_a = 16'b0000000000001101;
            14'h4e34: o_data_a = 16'b1110001100001000;
            14'h4e35: o_data_a = 16'b0100110110001010;
            14'h4e36: o_data_a = 16'b1110110000010000;
            14'h4e37: o_data_a = 16'b0000000000001110;
            14'h4e38: o_data_a = 16'b1110001100001000;
            14'h4e39: o_data_a = 16'b0100111000111101;
            14'h4e3a: o_data_a = 16'b1110110000010000;
            14'h4e3b: o_data_a = 16'b0000000001011111;
            14'h4e3c: o_data_a = 16'b1110101010000111;
            14'h4e3d: o_data_a = 16'b0000000000000000;
            14'h4e3e: o_data_a = 16'b1111110010101000;
            14'h4e3f: o_data_a = 16'b1111110000010000;
            14'h4e40: o_data_a = 16'b0000000000000101;
            14'h4e41: o_data_a = 16'b1110001100001000;
            14'h4e42: o_data_a = 16'b0000000000000000;
            14'h4e43: o_data_a = 16'b1111110111001000;
            14'h4e44: o_data_a = 16'b1111110010100000;
            14'h4e45: o_data_a = 16'b1110101010001000;
            14'h4e46: o_data_a = 16'b0000000000110110;
            14'h4e47: o_data_a = 16'b1110101010000111;
            14'h4e48: o_data_a = 16'b0000000000010110;
            14'h4e49: o_data_a = 16'b1111110000010000;
            14'h4e4a: o_data_a = 16'b0000000000000000;
            14'h4e4b: o_data_a = 16'b1111110111101000;
            14'h4e4c: o_data_a = 16'b1110110010100000;
            14'h4e4d: o_data_a = 16'b1110001100001000;
            14'h4e4e: o_data_a = 16'b0000000101100000;
            14'h4e4f: o_data_a = 16'b1110110000010000;
            14'h4e50: o_data_a = 16'b0000000000000000;
            14'h4e51: o_data_a = 16'b1111110111101000;
            14'h4e52: o_data_a = 16'b1110110010100000;
            14'h4e53: o_data_a = 16'b1110001100001000;
            14'h4e54: o_data_a = 16'b0000000000000000;
            14'h4e55: o_data_a = 16'b1111110010101000;
            14'h4e56: o_data_a = 16'b1111110000010000;
            14'h4e57: o_data_a = 16'b1110110010100000;
            14'h4e58: o_data_a = 16'b1111000010001000;
            14'h4e59: o_data_a = 16'b0000000000010111;
            14'h4e5a: o_data_a = 16'b1111110000010000;
            14'h4e5b: o_data_a = 16'b0000000000000000;
            14'h4e5c: o_data_a = 16'b1111110111101000;
            14'h4e5d: o_data_a = 16'b1110110010100000;
            14'h4e5e: o_data_a = 16'b1110001100001000;
            14'h4e5f: o_data_a = 16'b0000000000000000;
            14'h4e60: o_data_a = 16'b1111110010101000;
            14'h4e61: o_data_a = 16'b1111110000010000;
            14'h4e62: o_data_a = 16'b1110110010100000;
            14'h4e63: o_data_a = 16'b1111000111001000;
            14'h4e64: o_data_a = 16'b0000000000000000;
            14'h4e65: o_data_a = 16'b1111110010101000;
            14'h4e66: o_data_a = 16'b1111110000010000;
            14'h4e67: o_data_a = 16'b0000000000010110;
            14'h4e68: o_data_a = 16'b1110001100001000;
            14'h4e69: o_data_a = 16'b0000000000000000;
            14'h4e6a: o_data_a = 16'b1111110111001000;
            14'h4e6b: o_data_a = 16'b1111110010100000;
            14'h4e6c: o_data_a = 16'b1110101010001000;
            14'h4e6d: o_data_a = 16'b0000000000000000;
            14'h4e6e: o_data_a = 16'b1111110010101000;
            14'h4e6f: o_data_a = 16'b1111110000010000;
            14'h4e70: o_data_a = 16'b0000000000010111;
            14'h4e71: o_data_a = 16'b1110001100001000;
            14'h4e72: o_data_a = 16'b0000000000000000;
            14'h4e73: o_data_a = 16'b1111110111001000;
            14'h4e74: o_data_a = 16'b1111110010100000;
            14'h4e75: o_data_a = 16'b1110101010001000;
            14'h4e76: o_data_a = 16'b0000000000000000;
            14'h4e77: o_data_a = 16'b1111110010100000;
            14'h4e78: o_data_a = 16'b1111110001001000;
            14'h4e79: o_data_a = 16'b0000000000000000;
            14'h4e7a: o_data_a = 16'b1111110010101000;
            14'h4e7b: o_data_a = 16'b1111110000010000;
            14'h4e7c: o_data_a = 16'b0000000000010101;
            14'h4e7d: o_data_a = 16'b1110001100001000;
            14'h4e7e: o_data_a = 16'b0000000000010110;
            14'h4e7f: o_data_a = 16'b1111110000010000;
            14'h4e80: o_data_a = 16'b0000000000000000;
            14'h4e81: o_data_a = 16'b1111110111101000;
            14'h4e82: o_data_a = 16'b1110110010100000;
            14'h4e83: o_data_a = 16'b1110001100001000;
            14'h4e84: o_data_a = 16'b0001111111000000;
            14'h4e85: o_data_a = 16'b1110110000010000;
            14'h4e86: o_data_a = 16'b0000000000000000;
            14'h4e87: o_data_a = 16'b1111110111101000;
            14'h4e88: o_data_a = 16'b1110110010100000;
            14'h4e89: o_data_a = 16'b1110001100001000;
            14'h4e8a: o_data_a = 16'b0100111010001110;
            14'h4e8b: o_data_a = 16'b1110110000010000;
            14'h4e8c: o_data_a = 16'b0000000000000110;
            14'h4e8d: o_data_a = 16'b1110101010000111;
            14'h4e8e: o_data_a = 16'b0000000000000000;
            14'h4e8f: o_data_a = 16'b1111110010101000;
            14'h4e90: o_data_a = 16'b1111110000010000;
            14'h4e91: o_data_a = 16'b0100111010010101;
            14'h4e92: o_data_a = 16'b1110001100000101;
            14'h4e93: o_data_a = 16'b0100111010100000;
            14'h4e94: o_data_a = 16'b1110101010000111;
            14'h4e95: o_data_a = 16'b0000000000100000;
            14'h4e96: o_data_a = 16'b1110110000010000;
            14'h4e97: o_data_a = 16'b0000000000000000;
            14'h4e98: o_data_a = 16'b1111110111101000;
            14'h4e99: o_data_a = 16'b1110110010100000;
            14'h4e9a: o_data_a = 16'b1110001100001000;
            14'h4e9b: o_data_a = 16'b0000000000000000;
            14'h4e9c: o_data_a = 16'b1111110010101000;
            14'h4e9d: o_data_a = 16'b1111110000010000;
            14'h4e9e: o_data_a = 16'b0000000000010110;
            14'h4e9f: o_data_a = 16'b1110001100001000;
            14'h4ea0: o_data_a = 16'b0000000000000000;
            14'h4ea1: o_data_a = 16'b1111110111001000;
            14'h4ea2: o_data_a = 16'b1111110010100000;
            14'h4ea3: o_data_a = 16'b1110101010001000;
            14'h4ea4: o_data_a = 16'b0000000000110110;
            14'h4ea5: o_data_a = 16'b1110101010000111;
            14'h4ea6: o_data_a = 16'b0000000000010101;
            14'h4ea7: o_data_a = 16'b1111110000010000;
            14'h4ea8: o_data_a = 16'b0000000000000000;
            14'h4ea9: o_data_a = 16'b1111110111101000;
            14'h4eaa: o_data_a = 16'b1110110010100000;
            14'h4eab: o_data_a = 16'b1110001100001000;
            14'h4eac: o_data_a = 16'b0000000000000000;
            14'h4ead: o_data_a = 16'b1111110010101000;
            14'h4eae: o_data_a = 16'b1111110000010000;
            14'h4eaf: o_data_a = 16'b0100111010110011;
            14'h4eb0: o_data_a = 16'b1110001100000101;
            14'h4eb1: o_data_a = 16'b0100111101000000;
            14'h4eb2: o_data_a = 16'b1110101010000111;
            14'h4eb3: o_data_a = 16'b0000000000010111;
            14'h4eb4: o_data_a = 16'b1111110000010000;
            14'h4eb5: o_data_a = 16'b0000000000000000;
            14'h4eb6: o_data_a = 16'b1111110111101000;
            14'h4eb7: o_data_a = 16'b1110110010100000;
            14'h4eb8: o_data_a = 16'b1110001100001000;
            14'h4eb9: o_data_a = 16'b0000000000000000;
            14'h4eba: o_data_a = 16'b1111110111001000;
            14'h4ebb: o_data_a = 16'b1111110010100000;
            14'h4ebc: o_data_a = 16'b1110101010001000;
            14'h4ebd: o_data_a = 16'b0100111011000001;
            14'h4ebe: o_data_a = 16'b1110110000010000;
            14'h4ebf: o_data_a = 16'b0000000000010110;
            14'h4ec0: o_data_a = 16'b1110101010000111;
            14'h4ec1: o_data_a = 16'b0000000000000000;
            14'h4ec2: o_data_a = 16'b1111110010101000;
            14'h4ec3: o_data_a = 16'b1111110000010000;
            14'h4ec4: o_data_a = 16'b0100111011001000;
            14'h4ec5: o_data_a = 16'b1110001100000101;
            14'h4ec6: o_data_a = 16'b0100111011110010;
            14'h4ec7: o_data_a = 16'b1110101010000111;
            14'h4ec8: o_data_a = 16'b0000000000010111;
            14'h4ec9: o_data_a = 16'b1111110000010000;
            14'h4eca: o_data_a = 16'b0000000000000000;
            14'h4ecb: o_data_a = 16'b1111110111101000;
            14'h4ecc: o_data_a = 16'b1110110010100000;
            14'h4ecd: o_data_a = 16'b1110001100001000;
            14'h4ece: o_data_a = 16'b0000000000000000;
            14'h4ecf: o_data_a = 16'b1111110111001000;
            14'h4ed0: o_data_a = 16'b1111110010100000;
            14'h4ed1: o_data_a = 16'b1110111111001000;
            14'h4ed2: o_data_a = 16'b0000000000000000;
            14'h4ed3: o_data_a = 16'b1111110010101000;
            14'h4ed4: o_data_a = 16'b1111110000010000;
            14'h4ed5: o_data_a = 16'b1110110010100000;
            14'h4ed6: o_data_a = 16'b1111000111001000;
            14'h4ed7: o_data_a = 16'b0000000000000000;
            14'h4ed8: o_data_a = 16'b1111110010101000;
            14'h4ed9: o_data_a = 16'b1111110000010000;
            14'h4eda: o_data_a = 16'b0000000000010111;
            14'h4edb: o_data_a = 16'b1110001100001000;
            14'h4edc: o_data_a = 16'b0000000000010110;
            14'h4edd: o_data_a = 16'b1111110000010000;
            14'h4ede: o_data_a = 16'b0000000000000000;
            14'h4edf: o_data_a = 16'b1111110111101000;
            14'h4ee0: o_data_a = 16'b1110110010100000;
            14'h4ee1: o_data_a = 16'b1110001100001000;
            14'h4ee2: o_data_a = 16'b0000000000000000;
            14'h4ee3: o_data_a = 16'b1111110111001000;
            14'h4ee4: o_data_a = 16'b1111110010100000;
            14'h4ee5: o_data_a = 16'b1110111111001000;
            14'h4ee6: o_data_a = 16'b0000000000000000;
            14'h4ee7: o_data_a = 16'b1111110010101000;
            14'h4ee8: o_data_a = 16'b1111110000010000;
            14'h4ee9: o_data_a = 16'b1110110010100000;
            14'h4eea: o_data_a = 16'b1111000111001000;
            14'h4eeb: o_data_a = 16'b0000000000000000;
            14'h4eec: o_data_a = 16'b1111110010101000;
            14'h4eed: o_data_a = 16'b1111110000010000;
            14'h4eee: o_data_a = 16'b0000000000010110;
            14'h4eef: o_data_a = 16'b1110001100001000;
            14'h4ef0: o_data_a = 16'b0100111100110101;
            14'h4ef1: o_data_a = 16'b1110101010000111;
            14'h4ef2: o_data_a = 16'b0000000000011111;
            14'h4ef3: o_data_a = 16'b1110110000010000;
            14'h4ef4: o_data_a = 16'b0000000000000000;
            14'h4ef5: o_data_a = 16'b1111110111101000;
            14'h4ef6: o_data_a = 16'b1110110010100000;
            14'h4ef7: o_data_a = 16'b1110001100001000;
            14'h4ef8: o_data_a = 16'b0000000000000000;
            14'h4ef9: o_data_a = 16'b1111110010101000;
            14'h4efa: o_data_a = 16'b1111110000010000;
            14'h4efb: o_data_a = 16'b0000000000010111;
            14'h4efc: o_data_a = 16'b1110001100001000;
            14'h4efd: o_data_a = 16'b0000000000010110;
            14'h4efe: o_data_a = 16'b1111110000010000;
            14'h4eff: o_data_a = 16'b0000000000000000;
            14'h4f00: o_data_a = 16'b1111110111101000;
            14'h4f01: o_data_a = 16'b1110110010100000;
            14'h4f02: o_data_a = 16'b1110001100001000;
            14'h4f03: o_data_a = 16'b0000000000100000;
            14'h4f04: o_data_a = 16'b1110110000010000;
            14'h4f05: o_data_a = 16'b0000000000000000;
            14'h4f06: o_data_a = 16'b1111110111101000;
            14'h4f07: o_data_a = 16'b1110110010100000;
            14'h4f08: o_data_a = 16'b1110001100001000;
            14'h4f09: o_data_a = 16'b0100111100001101;
            14'h4f0a: o_data_a = 16'b1110110000010000;
            14'h4f0b: o_data_a = 16'b0000000000000110;
            14'h4f0c: o_data_a = 16'b1110101010000111;
            14'h4f0d: o_data_a = 16'b0000000000000000;
            14'h4f0e: o_data_a = 16'b1111110010101000;
            14'h4f0f: o_data_a = 16'b1111110000010000;
            14'h4f10: o_data_a = 16'b0100111100010100;
            14'h4f11: o_data_a = 16'b1110001100000101;
            14'h4f12: o_data_a = 16'b0100111100011111;
            14'h4f13: o_data_a = 16'b1110101010000111;
            14'h4f14: o_data_a = 16'b0001111111000000;
            14'h4f15: o_data_a = 16'b1110110000010000;
            14'h4f16: o_data_a = 16'b0000000000000000;
            14'h4f17: o_data_a = 16'b1111110111101000;
            14'h4f18: o_data_a = 16'b1110110010100000;
            14'h4f19: o_data_a = 16'b1110001100001000;
            14'h4f1a: o_data_a = 16'b0000000000000000;
            14'h4f1b: o_data_a = 16'b1111110010101000;
            14'h4f1c: o_data_a = 16'b1111110000010000;
            14'h4f1d: o_data_a = 16'b0000000000010110;
            14'h4f1e: o_data_a = 16'b1110001100001000;
            14'h4f1f: o_data_a = 16'b0000000000010110;
            14'h4f20: o_data_a = 16'b1111110000010000;
            14'h4f21: o_data_a = 16'b0000000000000000;
            14'h4f22: o_data_a = 16'b1111110111101000;
            14'h4f23: o_data_a = 16'b1110110010100000;
            14'h4f24: o_data_a = 16'b1110001100001000;
            14'h4f25: o_data_a = 16'b0000000101000001;
            14'h4f26: o_data_a = 16'b1110110000010000;
            14'h4f27: o_data_a = 16'b0000000000000000;
            14'h4f28: o_data_a = 16'b1111110111101000;
            14'h4f29: o_data_a = 16'b1110110010100000;
            14'h4f2a: o_data_a = 16'b1110001100001000;
            14'h4f2b: o_data_a = 16'b0000000000000000;
            14'h4f2c: o_data_a = 16'b1111110010101000;
            14'h4f2d: o_data_a = 16'b1111110000010000;
            14'h4f2e: o_data_a = 16'b1110110010100000;
            14'h4f2f: o_data_a = 16'b1111000111001000;
            14'h4f30: o_data_a = 16'b0000000000000000;
            14'h4f31: o_data_a = 16'b1111110010101000;
            14'h4f32: o_data_a = 16'b1111110000010000;
            14'h4f33: o_data_a = 16'b0000000000010110;
            14'h4f34: o_data_a = 16'b1110001100001000;
            14'h4f35: o_data_a = 16'b0000000000000000;
            14'h4f36: o_data_a = 16'b1111110111001000;
            14'h4f37: o_data_a = 16'b1111110010100000;
            14'h4f38: o_data_a = 16'b1110101010001000;
            14'h4f39: o_data_a = 16'b0000000000000000;
            14'h4f3a: o_data_a = 16'b1111110010101000;
            14'h4f3b: o_data_a = 16'b1111110000010000;
            14'h4f3c: o_data_a = 16'b0000000000010101;
            14'h4f3d: o_data_a = 16'b1110001100001000;
            14'h4f3e: o_data_a = 16'b0100111101001100;
            14'h4f3f: o_data_a = 16'b1110101010000111;
            14'h4f40: o_data_a = 16'b0000000000000000;
            14'h4f41: o_data_a = 16'b1111110111001000;
            14'h4f42: o_data_a = 16'b1111110010100000;
            14'h4f43: o_data_a = 16'b1110101010001000;
            14'h4f44: o_data_a = 16'b0000000000000000;
            14'h4f45: o_data_a = 16'b1111110010100000;
            14'h4f46: o_data_a = 16'b1111110001001000;
            14'h4f47: o_data_a = 16'b0000000000000000;
            14'h4f48: o_data_a = 16'b1111110010101000;
            14'h4f49: o_data_a = 16'b1111110000010000;
            14'h4f4a: o_data_a = 16'b0000000000010101;
            14'h4f4b: o_data_a = 16'b1110001100001000;
            14'h4f4c: o_data_a = 16'b0000000000100000;
            14'h4f4d: o_data_a = 16'b1110110000010000;
            14'h4f4e: o_data_a = 16'b0000000000000000;
            14'h4f4f: o_data_a = 16'b1111110111101000;
            14'h4f50: o_data_a = 16'b1110110010100000;
            14'h4f51: o_data_a = 16'b1110001100001000;
            14'h4f52: o_data_a = 16'b0000000000000001;
            14'h4f53: o_data_a = 16'b1110110000010000;
            14'h4f54: o_data_a = 16'b0000000000001101;
            14'h4f55: o_data_a = 16'b1110001100001000;
            14'h4f56: o_data_a = 16'b0100101001001101;
            14'h4f57: o_data_a = 16'b1110110000010000;
            14'h4f58: o_data_a = 16'b0000000000001110;
            14'h4f59: o_data_a = 16'b1110001100001000;
            14'h4f5a: o_data_a = 16'b0100111101011110;
            14'h4f5b: o_data_a = 16'b1110110000010000;
            14'h4f5c: o_data_a = 16'b0000000001011111;
            14'h4f5d: o_data_a = 16'b1110101010000111;
            14'h4f5e: o_data_a = 16'b0000000000000000;
            14'h4f5f: o_data_a = 16'b1111110010101000;
            14'h4f60: o_data_a = 16'b1111110000010000;
            14'h4f61: o_data_a = 16'b0000000000000101;
            14'h4f62: o_data_a = 16'b1110001100001000;
            14'h4f63: o_data_a = 16'b0000000000000000;
            14'h4f64: o_data_a = 16'b1111110111001000;
            14'h4f65: o_data_a = 16'b1111110010100000;
            14'h4f66: o_data_a = 16'b1110101010001000;
            14'h4f67: o_data_a = 16'b0000000000110110;
            14'h4f68: o_data_a = 16'b1110101010000111;
            14'h4f69: o_data_a = 16'b0000000000000000;
            14'h4f6a: o_data_a = 16'b1111110111101000;
            14'h4f6b: o_data_a = 16'b1110110010100000;
            14'h4f6c: o_data_a = 16'b1110101010001000;
            14'h4f6d: o_data_a = 16'b0100000000000000;
            14'h4f6e: o_data_a = 16'b1110110000010000;
            14'h4f6f: o_data_a = 16'b0000000000000000;
            14'h4f70: o_data_a = 16'b1111110111101000;
            14'h4f71: o_data_a = 16'b1110110010100000;
            14'h4f72: o_data_a = 16'b1110001100001000;
            14'h4f73: o_data_a = 16'b0000000000000000;
            14'h4f74: o_data_a = 16'b1111110010101000;
            14'h4f75: o_data_a = 16'b1111110000010000;
            14'h4f76: o_data_a = 16'b0000000000011011;
            14'h4f77: o_data_a = 16'b1110001100001000;
            14'h4f78: o_data_a = 16'b0000000000000000;
            14'h4f79: o_data_a = 16'b1111110111001000;
            14'h4f7a: o_data_a = 16'b1111110010100000;
            14'h4f7b: o_data_a = 16'b1110101010001000;
            14'h4f7c: o_data_a = 16'b0000000000000000;
            14'h4f7d: o_data_a = 16'b1111110010100000;
            14'h4f7e: o_data_a = 16'b1111110001001000;
            14'h4f7f: o_data_a = 16'b0000000000000000;
            14'h4f80: o_data_a = 16'b1111110010101000;
            14'h4f81: o_data_a = 16'b1111110000010000;
            14'h4f82: o_data_a = 16'b0000000000011100;
            14'h4f83: o_data_a = 16'b1110001100001000;
            14'h4f84: o_data_a = 16'b0000000000010001;
            14'h4f85: o_data_a = 16'b1110110000010000;
            14'h4f86: o_data_a = 16'b0000000000000000;
            14'h4f87: o_data_a = 16'b1111110111101000;
            14'h4f88: o_data_a = 16'b1110110010100000;
            14'h4f89: o_data_a = 16'b1110001100001000;
            14'h4f8a: o_data_a = 16'b0000000000000001;
            14'h4f8b: o_data_a = 16'b1110110000010000;
            14'h4f8c: o_data_a = 16'b0000000000001101;
            14'h4f8d: o_data_a = 16'b1110001100001000;
            14'h4f8e: o_data_a = 16'b0001011010110000;
            14'h4f8f: o_data_a = 16'b1110110000010000;
            14'h4f90: o_data_a = 16'b0000000000001110;
            14'h4f91: o_data_a = 16'b1110001100001000;
            14'h4f92: o_data_a = 16'b0100111110010110;
            14'h4f93: o_data_a = 16'b1110110000010000;
            14'h4f94: o_data_a = 16'b0000000001011111;
            14'h4f95: o_data_a = 16'b1110101010000111;
            14'h4f96: o_data_a = 16'b0000000000000000;
            14'h4f97: o_data_a = 16'b1111110010101000;
            14'h4f98: o_data_a = 16'b1111110000010000;
            14'h4f99: o_data_a = 16'b0000000000011101;
            14'h4f9a: o_data_a = 16'b1110001100001000;
            14'h4f9b: o_data_a = 16'b0000000000000000;
            14'h4f9c: o_data_a = 16'b1111110111001000;
            14'h4f9d: o_data_a = 16'b1111110010100000;
            14'h4f9e: o_data_a = 16'b1110101010001000;
            14'h4f9f: o_data_a = 16'b0000000000011101;
            14'h4fa0: o_data_a = 16'b1111110000010000;
            14'h4fa1: o_data_a = 16'b0000000000000000;
            14'h4fa2: o_data_a = 16'b1111110111101000;
            14'h4fa3: o_data_a = 16'b1110110010100000;
            14'h4fa4: o_data_a = 16'b1110001100001000;
            14'h4fa5: o_data_a = 16'b0000000000000000;
            14'h4fa6: o_data_a = 16'b1111110010101000;
            14'h4fa7: o_data_a = 16'b1111110000010000;
            14'h4fa8: o_data_a = 16'b1110110010100000;
            14'h4fa9: o_data_a = 16'b1111000010001000;
            14'h4faa: o_data_a = 16'b0000000000000000;
            14'h4fab: o_data_a = 16'b1111110111001000;
            14'h4fac: o_data_a = 16'b1111110010100000;
            14'h4fad: o_data_a = 16'b1110111111001000;
            14'h4fae: o_data_a = 16'b0000000000000000;
            14'h4faf: o_data_a = 16'b1111110010101000;
            14'h4fb0: o_data_a = 16'b1111110000010000;
            14'h4fb1: o_data_a = 16'b0000000000000101;
            14'h4fb2: o_data_a = 16'b1110001100001000;
            14'h4fb3: o_data_a = 16'b0000000000000000;
            14'h4fb4: o_data_a = 16'b1111110010101000;
            14'h4fb5: o_data_a = 16'b1111110000010000;
            14'h4fb6: o_data_a = 16'b0000000000000100;
            14'h4fb7: o_data_a = 16'b1110001100001000;
            14'h4fb8: o_data_a = 16'b0000000000000101;
            14'h4fb9: o_data_a = 16'b1111110000010000;
            14'h4fba: o_data_a = 16'b0000000000000000;
            14'h4fbb: o_data_a = 16'b1111110111101000;
            14'h4fbc: o_data_a = 16'b1110110010100000;
            14'h4fbd: o_data_a = 16'b1110001100001000;
            14'h4fbe: o_data_a = 16'b0000000000000000;
            14'h4fbf: o_data_a = 16'b1111110010101000;
            14'h4fc0: o_data_a = 16'b1111110000010000;
            14'h4fc1: o_data_a = 16'b0000000000000100;
            14'h4fc2: o_data_a = 16'b1111110000100000;
            14'h4fc3: o_data_a = 16'b1110001100001000;
            14'h4fc4: o_data_a = 16'b0000000000000001;
            14'h4fc5: o_data_a = 16'b1111110000100000;
            14'h4fc6: o_data_a = 16'b1111110000010000;
            14'h4fc7: o_data_a = 16'b0000000000000000;
            14'h4fc8: o_data_a = 16'b1111110111101000;
            14'h4fc9: o_data_a = 16'b1110110010100000;
            14'h4fca: o_data_a = 16'b1110001100001000;
            14'h4fcb: o_data_a = 16'b0000000000010000;
            14'h4fcc: o_data_a = 16'b1110110000010000;
            14'h4fcd: o_data_a = 16'b0000000000000000;
            14'h4fce: o_data_a = 16'b1111110111101000;
            14'h4fcf: o_data_a = 16'b1110110010100000;
            14'h4fd0: o_data_a = 16'b1110001100001000;
            14'h4fd1: o_data_a = 16'b0100111111010101;
            14'h4fd2: o_data_a = 16'b1110110000010000;
            14'h4fd3: o_data_a = 16'b0000000000100110;
            14'h4fd4: o_data_a = 16'b1110101010000111;
            14'h4fd5: o_data_a = 16'b0000000000000000;
            14'h4fd6: o_data_a = 16'b1111110010100000;
            14'h4fd7: o_data_a = 16'b1111110001001000;
            14'h4fd8: o_data_a = 16'b0000000000000000;
            14'h4fd9: o_data_a = 16'b1111110010101000;
            14'h4fda: o_data_a = 16'b1111110000010000;
            14'h4fdb: o_data_a = 16'b0101000001110000;
            14'h4fdc: o_data_a = 16'b1110001100000101;
            14'h4fdd: o_data_a = 16'b0000000000000001;
            14'h4fde: o_data_a = 16'b1111110000100000;
            14'h4fdf: o_data_a = 16'b1111110000010000;
            14'h4fe0: o_data_a = 16'b0000000000000000;
            14'h4fe1: o_data_a = 16'b1111110111101000;
            14'h4fe2: o_data_a = 16'b1110110010100000;
            14'h4fe3: o_data_a = 16'b1110001100001000;
            14'h4fe4: o_data_a = 16'b0000000000000000;
            14'h4fe5: o_data_a = 16'b1111110111001000;
            14'h4fe6: o_data_a = 16'b1111110010100000;
            14'h4fe7: o_data_a = 16'b1110111111001000;
            14'h4fe8: o_data_a = 16'b0000000000000000;
            14'h4fe9: o_data_a = 16'b1111110010101000;
            14'h4fea: o_data_a = 16'b1111110000010000;
            14'h4feb: o_data_a = 16'b1110110010100000;
            14'h4fec: o_data_a = 16'b1111000010001000;
            14'h4fed: o_data_a = 16'b0000000000000000;
            14'h4fee: o_data_a = 16'b1111110010101000;
            14'h4fef: o_data_a = 16'b1111110000010000;
            14'h4ff0: o_data_a = 16'b0000000000000001;
            14'h4ff1: o_data_a = 16'b1111110000100000;
            14'h4ff2: o_data_a = 16'b1110001100001000;
            14'h4ff3: o_data_a = 16'b0000000000000001;
            14'h4ff4: o_data_a = 16'b1111110000100000;
            14'h4ff5: o_data_a = 16'b1111110000010000;
            14'h4ff6: o_data_a = 16'b0000000000000000;
            14'h4ff7: o_data_a = 16'b1111110111101000;
            14'h4ff8: o_data_a = 16'b1110110010100000;
            14'h4ff9: o_data_a = 16'b1110001100001000;
            14'h4ffa: o_data_a = 16'b0000000000011101;
            14'h4ffb: o_data_a = 16'b1111110000010000;
            14'h4ffc: o_data_a = 16'b0000000000000000;
            14'h4ffd: o_data_a = 16'b1111110111101000;
            14'h4ffe: o_data_a = 16'b1110110010100000;
            14'h4fff: o_data_a = 16'b1110001100001000;
            14'h5000: o_data_a = 16'b0000000000000000;
            14'h5001: o_data_a = 16'b1111110010101000;
            14'h5002: o_data_a = 16'b1111110000010000;
            14'h5003: o_data_a = 16'b1110110010100000;
            14'h5004: o_data_a = 16'b1111000010001000;
            14'h5005: o_data_a = 16'b0000000000000001;
            14'h5006: o_data_a = 16'b1111110000100000;
            14'h5007: o_data_a = 16'b1111110000010000;
            14'h5008: o_data_a = 16'b0000000000000000;
            14'h5009: o_data_a = 16'b1111110111101000;
            14'h500a: o_data_a = 16'b1110110010100000;
            14'h500b: o_data_a = 16'b1110001100001000;
            14'h500c: o_data_a = 16'b0000000000000000;
            14'h500d: o_data_a = 16'b1111110111001000;
            14'h500e: o_data_a = 16'b1111110010100000;
            14'h500f: o_data_a = 16'b1110111111001000;
            14'h5010: o_data_a = 16'b0000000000000000;
            14'h5011: o_data_a = 16'b1111110010101000;
            14'h5012: o_data_a = 16'b1111110000010000;
            14'h5013: o_data_a = 16'b1110110010100000;
            14'h5014: o_data_a = 16'b1111000111001000;
            14'h5015: o_data_a = 16'b0000000000011101;
            14'h5016: o_data_a = 16'b1111110000010000;
            14'h5017: o_data_a = 16'b0000000000000000;
            14'h5018: o_data_a = 16'b1111110111101000;
            14'h5019: o_data_a = 16'b1110110010100000;
            14'h501a: o_data_a = 16'b1110001100001000;
            14'h501b: o_data_a = 16'b0000000000000000;
            14'h501c: o_data_a = 16'b1111110010101000;
            14'h501d: o_data_a = 16'b1111110000010000;
            14'h501e: o_data_a = 16'b1110110010100000;
            14'h501f: o_data_a = 16'b1111000010001000;
            14'h5020: o_data_a = 16'b0000000000000000;
            14'h5021: o_data_a = 16'b1111110010101000;
            14'h5022: o_data_a = 16'b1111110000010000;
            14'h5023: o_data_a = 16'b0000000000000100;
            14'h5024: o_data_a = 16'b1110001100001000;
            14'h5025: o_data_a = 16'b0000000000000100;
            14'h5026: o_data_a = 16'b1111110000100000;
            14'h5027: o_data_a = 16'b1111110000010000;
            14'h5028: o_data_a = 16'b0000000000000000;
            14'h5029: o_data_a = 16'b1111110111101000;
            14'h502a: o_data_a = 16'b1110110010100000;
            14'h502b: o_data_a = 16'b1110001100001000;
            14'h502c: o_data_a = 16'b0000000000000001;
            14'h502d: o_data_a = 16'b1111110000100000;
            14'h502e: o_data_a = 16'b1111110000010000;
            14'h502f: o_data_a = 16'b0000000000000000;
            14'h5030: o_data_a = 16'b1111110111101000;
            14'h5031: o_data_a = 16'b1110110010100000;
            14'h5032: o_data_a = 16'b1110001100001000;
            14'h5033: o_data_a = 16'b0000000000000000;
            14'h5034: o_data_a = 16'b1111110111001000;
            14'h5035: o_data_a = 16'b1111110010100000;
            14'h5036: o_data_a = 16'b1110111111001000;
            14'h5037: o_data_a = 16'b0000000000000000;
            14'h5038: o_data_a = 16'b1111110010101000;
            14'h5039: o_data_a = 16'b1111110000010000;
            14'h503a: o_data_a = 16'b1110110010100000;
            14'h503b: o_data_a = 16'b1111000111001000;
            14'h503c: o_data_a = 16'b0000000000011101;
            14'h503d: o_data_a = 16'b1111110000010000;
            14'h503e: o_data_a = 16'b0000000000000000;
            14'h503f: o_data_a = 16'b1111110111101000;
            14'h5040: o_data_a = 16'b1110110010100000;
            14'h5041: o_data_a = 16'b1110001100001000;
            14'h5042: o_data_a = 16'b0000000000000000;
            14'h5043: o_data_a = 16'b1111110010101000;
            14'h5044: o_data_a = 16'b1111110000010000;
            14'h5045: o_data_a = 16'b1110110010100000;
            14'h5046: o_data_a = 16'b1111000010001000;
            14'h5047: o_data_a = 16'b0000000000000000;
            14'h5048: o_data_a = 16'b1111110010101000;
            14'h5049: o_data_a = 16'b1111110000010000;
            14'h504a: o_data_a = 16'b0000000000000100;
            14'h504b: o_data_a = 16'b1110001100001000;
            14'h504c: o_data_a = 16'b0000000000000100;
            14'h504d: o_data_a = 16'b1111110000100000;
            14'h504e: o_data_a = 16'b1111110000010000;
            14'h504f: o_data_a = 16'b0000000000000000;
            14'h5050: o_data_a = 16'b1111110111101000;
            14'h5051: o_data_a = 16'b1110110010100000;
            14'h5052: o_data_a = 16'b1110001100001000;
            14'h5053: o_data_a = 16'b0000000000000000;
            14'h5054: o_data_a = 16'b1111110010101000;
            14'h5055: o_data_a = 16'b1111110000010000;
            14'h5056: o_data_a = 16'b1110110010100000;
            14'h5057: o_data_a = 16'b1111000010001000;
            14'h5058: o_data_a = 16'b0000000000000000;
            14'h5059: o_data_a = 16'b1111110010101000;
            14'h505a: o_data_a = 16'b1111110000010000;
            14'h505b: o_data_a = 16'b0000000000000101;
            14'h505c: o_data_a = 16'b1110001100001000;
            14'h505d: o_data_a = 16'b0000000000000000;
            14'h505e: o_data_a = 16'b1111110010101000;
            14'h505f: o_data_a = 16'b1111110000010000;
            14'h5060: o_data_a = 16'b0000000000000100;
            14'h5061: o_data_a = 16'b1110001100001000;
            14'h5062: o_data_a = 16'b0000000000000101;
            14'h5063: o_data_a = 16'b1111110000010000;
            14'h5064: o_data_a = 16'b0000000000000000;
            14'h5065: o_data_a = 16'b1111110111101000;
            14'h5066: o_data_a = 16'b1110110010100000;
            14'h5067: o_data_a = 16'b1110001100001000;
            14'h5068: o_data_a = 16'b0000000000000000;
            14'h5069: o_data_a = 16'b1111110010101000;
            14'h506a: o_data_a = 16'b1111110000010000;
            14'h506b: o_data_a = 16'b0000000000000100;
            14'h506c: o_data_a = 16'b1111110000100000;
            14'h506d: o_data_a = 16'b1110001100001000;
            14'h506e: o_data_a = 16'b0100111111000100;
            14'h506f: o_data_a = 16'b1110101010000111;
            14'h5070: o_data_a = 16'b0000000000000000;
            14'h5071: o_data_a = 16'b1111110111001000;
            14'h5072: o_data_a = 16'b1111110010100000;
            14'h5073: o_data_a = 16'b1110101010001000;
            14'h5074: o_data_a = 16'b0000000000110110;
            14'h5075: o_data_a = 16'b1110101010000111;
            14'h5076: o_data_a = 16'b0000000000000000;
            14'h5077: o_data_a = 16'b1111110111101000;
            14'h5078: o_data_a = 16'b1110110010100000;
            14'h5079: o_data_a = 16'b1110101010001000;
            14'h507a: o_data_a = 16'b0000000000000001;
            14'h507b: o_data_a = 16'b1111110000100000;
            14'h507c: o_data_a = 16'b1111110000010000;
            14'h507d: o_data_a = 16'b0000000000000000;
            14'h507e: o_data_a = 16'b1111110111101000;
            14'h507f: o_data_a = 16'b1110110010100000;
            14'h5080: o_data_a = 16'b1110001100001000;
            14'h5081: o_data_a = 16'b0010000000000000;
            14'h5082: o_data_a = 16'b1110110000010000;
            14'h5083: o_data_a = 16'b0000000000000000;
            14'h5084: o_data_a = 16'b1111110111101000;
            14'h5085: o_data_a = 16'b1110110010100000;
            14'h5086: o_data_a = 16'b1110001100001000;
            14'h5087: o_data_a = 16'b0101000010001011;
            14'h5088: o_data_a = 16'b1110110000010000;
            14'h5089: o_data_a = 16'b0000000000100110;
            14'h508a: o_data_a = 16'b1110101010000111;
            14'h508b: o_data_a = 16'b0000000000000000;
            14'h508c: o_data_a = 16'b1111110010100000;
            14'h508d: o_data_a = 16'b1111110001001000;
            14'h508e: o_data_a = 16'b0000000000000000;
            14'h508f: o_data_a = 16'b1111110010101000;
            14'h5090: o_data_a = 16'b1111110000010000;
            14'h5091: o_data_a = 16'b0101000011010111;
            14'h5092: o_data_a = 16'b1110001100000101;
            14'h5093: o_data_a = 16'b0000000000000001;
            14'h5094: o_data_a = 16'b1111110000100000;
            14'h5095: o_data_a = 16'b1111110000010000;
            14'h5096: o_data_a = 16'b0000000000000000;
            14'h5097: o_data_a = 16'b1111110111101000;
            14'h5098: o_data_a = 16'b1110110010100000;
            14'h5099: o_data_a = 16'b1110001100001000;
            14'h509a: o_data_a = 16'b0000000000011011;
            14'h509b: o_data_a = 16'b1111110000010000;
            14'h509c: o_data_a = 16'b0000000000000000;
            14'h509d: o_data_a = 16'b1111110111101000;
            14'h509e: o_data_a = 16'b1110110010100000;
            14'h509f: o_data_a = 16'b1110001100001000;
            14'h50a0: o_data_a = 16'b0000000000000000;
            14'h50a1: o_data_a = 16'b1111110010101000;
            14'h50a2: o_data_a = 16'b1111110000010000;
            14'h50a3: o_data_a = 16'b1110110010100000;
            14'h50a4: o_data_a = 16'b1111000010001000;
            14'h50a5: o_data_a = 16'b0000000000000000;
            14'h50a6: o_data_a = 16'b1111110111001000;
            14'h50a7: o_data_a = 16'b1111110010100000;
            14'h50a8: o_data_a = 16'b1110101010001000;
            14'h50a9: o_data_a = 16'b0000000000000000;
            14'h50aa: o_data_a = 16'b1111110010101000;
            14'h50ab: o_data_a = 16'b1111110000010000;
            14'h50ac: o_data_a = 16'b0000000000000101;
            14'h50ad: o_data_a = 16'b1110001100001000;
            14'h50ae: o_data_a = 16'b0000000000000000;
            14'h50af: o_data_a = 16'b1111110010101000;
            14'h50b0: o_data_a = 16'b1111110000010000;
            14'h50b1: o_data_a = 16'b0000000000000100;
            14'h50b2: o_data_a = 16'b1110001100001000;
            14'h50b3: o_data_a = 16'b0000000000000101;
            14'h50b4: o_data_a = 16'b1111110000010000;
            14'h50b5: o_data_a = 16'b0000000000000000;
            14'h50b6: o_data_a = 16'b1111110111101000;
            14'h50b7: o_data_a = 16'b1110110010100000;
            14'h50b8: o_data_a = 16'b1110001100001000;
            14'h50b9: o_data_a = 16'b0000000000000000;
            14'h50ba: o_data_a = 16'b1111110010101000;
            14'h50bb: o_data_a = 16'b1111110000010000;
            14'h50bc: o_data_a = 16'b0000000000000100;
            14'h50bd: o_data_a = 16'b1111110000100000;
            14'h50be: o_data_a = 16'b1110001100001000;
            14'h50bf: o_data_a = 16'b0000000000000001;
            14'h50c0: o_data_a = 16'b1111110000100000;
            14'h50c1: o_data_a = 16'b1111110000010000;
            14'h50c2: o_data_a = 16'b0000000000000000;
            14'h50c3: o_data_a = 16'b1111110111101000;
            14'h50c4: o_data_a = 16'b1110110010100000;
            14'h50c5: o_data_a = 16'b1110001100001000;
            14'h50c6: o_data_a = 16'b0000000000000000;
            14'h50c7: o_data_a = 16'b1111110111001000;
            14'h50c8: o_data_a = 16'b1111110010100000;
            14'h50c9: o_data_a = 16'b1110111111001000;
            14'h50ca: o_data_a = 16'b0000000000000000;
            14'h50cb: o_data_a = 16'b1111110010101000;
            14'h50cc: o_data_a = 16'b1111110000010000;
            14'h50cd: o_data_a = 16'b1110110010100000;
            14'h50ce: o_data_a = 16'b1111000010001000;
            14'h50cf: o_data_a = 16'b0000000000000000;
            14'h50d0: o_data_a = 16'b1111110010101000;
            14'h50d1: o_data_a = 16'b1111110000010000;
            14'h50d2: o_data_a = 16'b0000000000000001;
            14'h50d3: o_data_a = 16'b1111110000100000;
            14'h50d4: o_data_a = 16'b1110001100001000;
            14'h50d5: o_data_a = 16'b0101000001111010;
            14'h50d6: o_data_a = 16'b1110101010000111;
            14'h50d7: o_data_a = 16'b0000000000000000;
            14'h50d8: o_data_a = 16'b1111110111001000;
            14'h50d9: o_data_a = 16'b1111110010100000;
            14'h50da: o_data_a = 16'b1110101010001000;
            14'h50db: o_data_a = 16'b0000000000110110;
            14'h50dc: o_data_a = 16'b1110101010000111;
            14'h50dd: o_data_a = 16'b0000000000011100;
            14'h50de: o_data_a = 16'b1111110000010000;
            14'h50df: o_data_a = 16'b0000000000000000;
            14'h50e0: o_data_a = 16'b1111110111101000;
            14'h50e1: o_data_a = 16'b1110110010100000;
            14'h50e2: o_data_a = 16'b1110001100001000;
            14'h50e3: o_data_a = 16'b0000000000000000;
            14'h50e4: o_data_a = 16'b1111110010101000;
            14'h50e5: o_data_a = 16'b1111110000010000;
            14'h50e6: o_data_a = 16'b0101000011101010;
            14'h50e7: o_data_a = 16'b1110001100000101;
            14'h50e8: o_data_a = 16'b0101000100111110;
            14'h50e9: o_data_a = 16'b1110101010000111;
            14'h50ea: o_data_a = 16'b0000000000000010;
            14'h50eb: o_data_a = 16'b1111110000100000;
            14'h50ec: o_data_a = 16'b1111110000010000;
            14'h50ed: o_data_a = 16'b0000000000000000;
            14'h50ee: o_data_a = 16'b1111110111101000;
            14'h50ef: o_data_a = 16'b1110110010100000;
            14'h50f0: o_data_a = 16'b1110001100001000;
            14'h50f1: o_data_a = 16'b0000000000011011;
            14'h50f2: o_data_a = 16'b1111110000010000;
            14'h50f3: o_data_a = 16'b0000000000000000;
            14'h50f4: o_data_a = 16'b1111110111101000;
            14'h50f5: o_data_a = 16'b1110110010100000;
            14'h50f6: o_data_a = 16'b1110001100001000;
            14'h50f7: o_data_a = 16'b0000000000000000;
            14'h50f8: o_data_a = 16'b1111110010101000;
            14'h50f9: o_data_a = 16'b1111110000010000;
            14'h50fa: o_data_a = 16'b1110110010100000;
            14'h50fb: o_data_a = 16'b1111000010001000;
            14'h50fc: o_data_a = 16'b0000000000000010;
            14'h50fd: o_data_a = 16'b1111110000100000;
            14'h50fe: o_data_a = 16'b1111110000010000;
            14'h50ff: o_data_a = 16'b0000000000000000;
            14'h5100: o_data_a = 16'b1111110111101000;
            14'h5101: o_data_a = 16'b1110110010100000;
            14'h5102: o_data_a = 16'b1110001100001000;
            14'h5103: o_data_a = 16'b0000000000011011;
            14'h5104: o_data_a = 16'b1111110000010000;
            14'h5105: o_data_a = 16'b0000000000000000;
            14'h5106: o_data_a = 16'b1111110111101000;
            14'h5107: o_data_a = 16'b1110110010100000;
            14'h5108: o_data_a = 16'b1110001100001000;
            14'h5109: o_data_a = 16'b0000000000000000;
            14'h510a: o_data_a = 16'b1111110010101000;
            14'h510b: o_data_a = 16'b1111110000010000;
            14'h510c: o_data_a = 16'b1110110010100000;
            14'h510d: o_data_a = 16'b1111000010001000;
            14'h510e: o_data_a = 16'b0000000000000000;
            14'h510f: o_data_a = 16'b1111110010101000;
            14'h5110: o_data_a = 16'b1111110000010000;
            14'h5111: o_data_a = 16'b0000000000000100;
            14'h5112: o_data_a = 16'b1110001100001000;
            14'h5113: o_data_a = 16'b0000000000000100;
            14'h5114: o_data_a = 16'b1111110000100000;
            14'h5115: o_data_a = 16'b1111110000010000;
            14'h5116: o_data_a = 16'b0000000000000000;
            14'h5117: o_data_a = 16'b1111110111101000;
            14'h5118: o_data_a = 16'b1110110010100000;
            14'h5119: o_data_a = 16'b1110001100001000;
            14'h511a: o_data_a = 16'b0000000000000010;
            14'h511b: o_data_a = 16'b1111110111100000;
            14'h511c: o_data_a = 16'b1111110000010000;
            14'h511d: o_data_a = 16'b0000000000000000;
            14'h511e: o_data_a = 16'b1111110111101000;
            14'h511f: o_data_a = 16'b1110110010100000;
            14'h5120: o_data_a = 16'b1110001100001000;
            14'h5121: o_data_a = 16'b0000000000000000;
            14'h5122: o_data_a = 16'b1111110010101000;
            14'h5123: o_data_a = 16'b1111110000010000;
            14'h5124: o_data_a = 16'b1110110010100000;
            14'h5125: o_data_a = 16'b1111010101001000;
            14'h5126: o_data_a = 16'b0000000000000000;
            14'h5127: o_data_a = 16'b1111110010101000;
            14'h5128: o_data_a = 16'b1111110000010000;
            14'h5129: o_data_a = 16'b0000000000000101;
            14'h512a: o_data_a = 16'b1110001100001000;
            14'h512b: o_data_a = 16'b0000000000000000;
            14'h512c: o_data_a = 16'b1111110010101000;
            14'h512d: o_data_a = 16'b1111110000010000;
            14'h512e: o_data_a = 16'b0000000000000100;
            14'h512f: o_data_a = 16'b1110001100001000;
            14'h5130: o_data_a = 16'b0000000000000101;
            14'h5131: o_data_a = 16'b1111110000010000;
            14'h5132: o_data_a = 16'b0000000000000000;
            14'h5133: o_data_a = 16'b1111110111101000;
            14'h5134: o_data_a = 16'b1110110010100000;
            14'h5135: o_data_a = 16'b1110001100001000;
            14'h5136: o_data_a = 16'b0000000000000000;
            14'h5137: o_data_a = 16'b1111110010101000;
            14'h5138: o_data_a = 16'b1111110000010000;
            14'h5139: o_data_a = 16'b0000000000000100;
            14'h513a: o_data_a = 16'b1111110000100000;
            14'h513b: o_data_a = 16'b1110001100001000;
            14'h513c: o_data_a = 16'b0101000110010011;
            14'h513d: o_data_a = 16'b1110101010000111;
            14'h513e: o_data_a = 16'b0000000000000010;
            14'h513f: o_data_a = 16'b1111110000100000;
            14'h5140: o_data_a = 16'b1111110000010000;
            14'h5141: o_data_a = 16'b0000000000000000;
            14'h5142: o_data_a = 16'b1111110111101000;
            14'h5143: o_data_a = 16'b1110110010100000;
            14'h5144: o_data_a = 16'b1110001100001000;
            14'h5145: o_data_a = 16'b0000000000011011;
            14'h5146: o_data_a = 16'b1111110000010000;
            14'h5147: o_data_a = 16'b0000000000000000;
            14'h5148: o_data_a = 16'b1111110111101000;
            14'h5149: o_data_a = 16'b1110110010100000;
            14'h514a: o_data_a = 16'b1110001100001000;
            14'h514b: o_data_a = 16'b0000000000000000;
            14'h514c: o_data_a = 16'b1111110010101000;
            14'h514d: o_data_a = 16'b1111110000010000;
            14'h514e: o_data_a = 16'b1110110010100000;
            14'h514f: o_data_a = 16'b1111000010001000;
            14'h5150: o_data_a = 16'b0000000000000010;
            14'h5151: o_data_a = 16'b1111110000100000;
            14'h5152: o_data_a = 16'b1111110000010000;
            14'h5153: o_data_a = 16'b0000000000000000;
            14'h5154: o_data_a = 16'b1111110111101000;
            14'h5155: o_data_a = 16'b1110110010100000;
            14'h5156: o_data_a = 16'b1110001100001000;
            14'h5157: o_data_a = 16'b0000000000011011;
            14'h5158: o_data_a = 16'b1111110000010000;
            14'h5159: o_data_a = 16'b0000000000000000;
            14'h515a: o_data_a = 16'b1111110111101000;
            14'h515b: o_data_a = 16'b1110110010100000;
            14'h515c: o_data_a = 16'b1110001100001000;
            14'h515d: o_data_a = 16'b0000000000000000;
            14'h515e: o_data_a = 16'b1111110010101000;
            14'h515f: o_data_a = 16'b1111110000010000;
            14'h5160: o_data_a = 16'b1110110010100000;
            14'h5161: o_data_a = 16'b1111000010001000;
            14'h5162: o_data_a = 16'b0000000000000000;
            14'h5163: o_data_a = 16'b1111110010101000;
            14'h5164: o_data_a = 16'b1111110000010000;
            14'h5165: o_data_a = 16'b0000000000000100;
            14'h5166: o_data_a = 16'b1110001100001000;
            14'h5167: o_data_a = 16'b0000000000000100;
            14'h5168: o_data_a = 16'b1111110000100000;
            14'h5169: o_data_a = 16'b1111110000010000;
            14'h516a: o_data_a = 16'b0000000000000000;
            14'h516b: o_data_a = 16'b1111110111101000;
            14'h516c: o_data_a = 16'b1110110010100000;
            14'h516d: o_data_a = 16'b1110001100001000;
            14'h516e: o_data_a = 16'b0000000000000010;
            14'h516f: o_data_a = 16'b1111110111100000;
            14'h5170: o_data_a = 16'b1111110000010000;
            14'h5171: o_data_a = 16'b0000000000000000;
            14'h5172: o_data_a = 16'b1111110111101000;
            14'h5173: o_data_a = 16'b1110110010100000;
            14'h5174: o_data_a = 16'b1110001100001000;
            14'h5175: o_data_a = 16'b0000000000000000;
            14'h5176: o_data_a = 16'b1111110010100000;
            14'h5177: o_data_a = 16'b1111110001001000;
            14'h5178: o_data_a = 16'b0000000000000000;
            14'h5179: o_data_a = 16'b1111110010101000;
            14'h517a: o_data_a = 16'b1111110000010000;
            14'h517b: o_data_a = 16'b1110110010100000;
            14'h517c: o_data_a = 16'b1111000000001000;
            14'h517d: o_data_a = 16'b0000000000000000;
            14'h517e: o_data_a = 16'b1111110010101000;
            14'h517f: o_data_a = 16'b1111110000010000;
            14'h5180: o_data_a = 16'b0000000000000101;
            14'h5181: o_data_a = 16'b1110001100001000;
            14'h5182: o_data_a = 16'b0000000000000000;
            14'h5183: o_data_a = 16'b1111110010101000;
            14'h5184: o_data_a = 16'b1111110000010000;
            14'h5185: o_data_a = 16'b0000000000000100;
            14'h5186: o_data_a = 16'b1110001100001000;
            14'h5187: o_data_a = 16'b0000000000000101;
            14'h5188: o_data_a = 16'b1111110000010000;
            14'h5189: o_data_a = 16'b0000000000000000;
            14'h518a: o_data_a = 16'b1111110111101000;
            14'h518b: o_data_a = 16'b1110110010100000;
            14'h518c: o_data_a = 16'b1110001100001000;
            14'h518d: o_data_a = 16'b0000000000000000;
            14'h518e: o_data_a = 16'b1111110010101000;
            14'h518f: o_data_a = 16'b1111110000010000;
            14'h5190: o_data_a = 16'b0000000000000100;
            14'h5191: o_data_a = 16'b1111110000100000;
            14'h5192: o_data_a = 16'b1110001100001000;
            14'h5193: o_data_a = 16'b0000000000000000;
            14'h5194: o_data_a = 16'b1111110111001000;
            14'h5195: o_data_a = 16'b1111110010100000;
            14'h5196: o_data_a = 16'b1110101010001000;
            14'h5197: o_data_a = 16'b0000000000110110;
            14'h5198: o_data_a = 16'b1110101010000111;
            14'h5199: o_data_a = 16'b0000000000000010;
            14'h519a: o_data_a = 16'b1111110000100000;
            14'h519b: o_data_a = 16'b1111110000010000;
            14'h519c: o_data_a = 16'b0000000000000000;
            14'h519d: o_data_a = 16'b1111110111101000;
            14'h519e: o_data_a = 16'b1110110010100000;
            14'h519f: o_data_a = 16'b1110001100001000;
            14'h51a0: o_data_a = 16'b0000000000000000;
            14'h51a1: o_data_a = 16'b1111110010101000;
            14'h51a2: o_data_a = 16'b1111110000010000;
            14'h51a3: o_data_a = 16'b0000000000011100;
            14'h51a4: o_data_a = 16'b1110001100001000;
            14'h51a5: o_data_a = 16'b0000000000000000;
            14'h51a6: o_data_a = 16'b1111110111001000;
            14'h51a7: o_data_a = 16'b1111110010100000;
            14'h51a8: o_data_a = 16'b1110101010001000;
            14'h51a9: o_data_a = 16'b0000000000110110;
            14'h51aa: o_data_a = 16'b1110101010000111;
            14'h51ab: o_data_a = 16'b0000000000000011;
            14'h51ac: o_data_a = 16'b1110110000010000;
            14'h51ad: o_data_a = 16'b1110001110010000;
            14'h51ae: o_data_a = 16'b0000000000000000;
            14'h51af: o_data_a = 16'b1111110111101000;
            14'h51b0: o_data_a = 16'b1110110010100000;
            14'h51b1: o_data_a = 16'b1110101010001000;
            14'h51b2: o_data_a = 16'b0101000110101101;
            14'h51b3: o_data_a = 16'b1110001100000001;
            14'h51b4: o_data_a = 16'b0000000000000010;
            14'h51b5: o_data_a = 16'b1111110000100000;
            14'h51b6: o_data_a = 16'b1111110000010000;
            14'h51b7: o_data_a = 16'b0000000000000000;
            14'h51b8: o_data_a = 16'b1111110111101000;
            14'h51b9: o_data_a = 16'b1110110010100000;
            14'h51ba: o_data_a = 16'b1110001100001000;
            14'h51bb: o_data_a = 16'b0000000000000000;
            14'h51bc: o_data_a = 16'b1111110111001000;
            14'h51bd: o_data_a = 16'b1111110010100000;
            14'h51be: o_data_a = 16'b1110101010001000;
            14'h51bf: o_data_a = 16'b0101000111000011;
            14'h51c0: o_data_a = 16'b1110110000010000;
            14'h51c1: o_data_a = 16'b0000000000100110;
            14'h51c2: o_data_a = 16'b1110101010000111;
            14'h51c3: o_data_a = 16'b0000000000000010;
            14'h51c4: o_data_a = 16'b1111110000100000;
            14'h51c5: o_data_a = 16'b1111110000010000;
            14'h51c6: o_data_a = 16'b0000000000000000;
            14'h51c7: o_data_a = 16'b1111110111101000;
            14'h51c8: o_data_a = 16'b1110110010100000;
            14'h51c9: o_data_a = 16'b1110001100001000;
            14'h51ca: o_data_a = 16'b0000000111111111;
            14'h51cb: o_data_a = 16'b1110110000010000;
            14'h51cc: o_data_a = 16'b0000000000000000;
            14'h51cd: o_data_a = 16'b1111110111101000;
            14'h51ce: o_data_a = 16'b1110110010100000;
            14'h51cf: o_data_a = 16'b1110001100001000;
            14'h51d0: o_data_a = 16'b0101000111010100;
            14'h51d1: o_data_a = 16'b1110110000010000;
            14'h51d2: o_data_a = 16'b0000000000010110;
            14'h51d3: o_data_a = 16'b1110101010000111;
            14'h51d4: o_data_a = 16'b0000000000000000;
            14'h51d5: o_data_a = 16'b1111110010101000;
            14'h51d6: o_data_a = 16'b1111110000010000;
            14'h51d7: o_data_a = 16'b1110110010100000;
            14'h51d8: o_data_a = 16'b1111010101001000;
            14'h51d9: o_data_a = 16'b0000000000000010;
            14'h51da: o_data_a = 16'b1111110111100000;
            14'h51db: o_data_a = 16'b1111110000010000;
            14'h51dc: o_data_a = 16'b0000000000000000;
            14'h51dd: o_data_a = 16'b1111110111101000;
            14'h51de: o_data_a = 16'b1110110010100000;
            14'h51df: o_data_a = 16'b1110001100001000;
            14'h51e0: o_data_a = 16'b0000000000000000;
            14'h51e1: o_data_a = 16'b1111110111001000;
            14'h51e2: o_data_a = 16'b1111110010100000;
            14'h51e3: o_data_a = 16'b1110101010001000;
            14'h51e4: o_data_a = 16'b0101000111101000;
            14'h51e5: o_data_a = 16'b1110110000010000;
            14'h51e6: o_data_a = 16'b0000000000100110;
            14'h51e7: o_data_a = 16'b1110101010000111;
            14'h51e8: o_data_a = 16'b0000000000000000;
            14'h51e9: o_data_a = 16'b1111110010101000;
            14'h51ea: o_data_a = 16'b1111110000010000;
            14'h51eb: o_data_a = 16'b1110110010100000;
            14'h51ec: o_data_a = 16'b1111010101001000;
            14'h51ed: o_data_a = 16'b0000000000000010;
            14'h51ee: o_data_a = 16'b1111110111100000;
            14'h51ef: o_data_a = 16'b1111110000010000;
            14'h51f0: o_data_a = 16'b0000000000000000;
            14'h51f1: o_data_a = 16'b1111110111101000;
            14'h51f2: o_data_a = 16'b1110110010100000;
            14'h51f3: o_data_a = 16'b1110001100001000;
            14'h51f4: o_data_a = 16'b0000000011111111;
            14'h51f5: o_data_a = 16'b1110110000010000;
            14'h51f6: o_data_a = 16'b0000000000000000;
            14'h51f7: o_data_a = 16'b1111110111101000;
            14'h51f8: o_data_a = 16'b1110110010100000;
            14'h51f9: o_data_a = 16'b1110001100001000;
            14'h51fa: o_data_a = 16'b0101000111111110;
            14'h51fb: o_data_a = 16'b1110110000010000;
            14'h51fc: o_data_a = 16'b0000000000010110;
            14'h51fd: o_data_a = 16'b1110101010000111;
            14'h51fe: o_data_a = 16'b0000000000000000;
            14'h51ff: o_data_a = 16'b1111110010101000;
            14'h5200: o_data_a = 16'b1111110000010000;
            14'h5201: o_data_a = 16'b1110110010100000;
            14'h5202: o_data_a = 16'b1111010101001000;
            14'h5203: o_data_a = 16'b0000000000000000;
            14'h5204: o_data_a = 16'b1111110010101000;
            14'h5205: o_data_a = 16'b1111110000010000;
            14'h5206: o_data_a = 16'b0101001000001010;
            14'h5207: o_data_a = 16'b1110001100000101;
            14'h5208: o_data_a = 16'b0101001000100001;
            14'h5209: o_data_a = 16'b1110101010000111;
            14'h520a: o_data_a = 16'b0000000000000111;
            14'h520b: o_data_a = 16'b1110110000010000;
            14'h520c: o_data_a = 16'b0000000000000000;
            14'h520d: o_data_a = 16'b1111110111101000;
            14'h520e: o_data_a = 16'b1110110010100000;
            14'h520f: o_data_a = 16'b1110001100001000;
            14'h5210: o_data_a = 16'b0000000000000001;
            14'h5211: o_data_a = 16'b1110110000010000;
            14'h5212: o_data_a = 16'b0000000000001101;
            14'h5213: o_data_a = 16'b1110001100001000;
            14'h5214: o_data_a = 16'b0110101011011001;
            14'h5215: o_data_a = 16'b1110110000010000;
            14'h5216: o_data_a = 16'b0000000000001110;
            14'h5217: o_data_a = 16'b1110001100001000;
            14'h5218: o_data_a = 16'b0101001000011100;
            14'h5219: o_data_a = 16'b1110110000010000;
            14'h521a: o_data_a = 16'b0000000001011111;
            14'h521b: o_data_a = 16'b1110101010000111;
            14'h521c: o_data_a = 16'b0000000000000000;
            14'h521d: o_data_a = 16'b1111110010101000;
            14'h521e: o_data_a = 16'b1111110000010000;
            14'h521f: o_data_a = 16'b0000000000000101;
            14'h5220: o_data_a = 16'b1110001100001000;
            14'h5221: o_data_a = 16'b0000000000000010;
            14'h5222: o_data_a = 16'b1111110000100000;
            14'h5223: o_data_a = 16'b1111110000010000;
            14'h5224: o_data_a = 16'b0000000000000000;
            14'h5225: o_data_a = 16'b1111110111101000;
            14'h5226: o_data_a = 16'b1110110010100000;
            14'h5227: o_data_a = 16'b1110001100001000;
            14'h5228: o_data_a = 16'b0000000000010000;
            14'h5229: o_data_a = 16'b1110110000010000;
            14'h522a: o_data_a = 16'b0000000000000000;
            14'h522b: o_data_a = 16'b1111110111101000;
            14'h522c: o_data_a = 16'b1110110010100000;
            14'h522d: o_data_a = 16'b1110001100001000;
            14'h522e: o_data_a = 16'b0000000000000010;
            14'h522f: o_data_a = 16'b1110110000010000;
            14'h5230: o_data_a = 16'b0000000000001101;
            14'h5231: o_data_a = 16'b1110001100001000;
            14'h5232: o_data_a = 16'b0001110001110111;
            14'h5233: o_data_a = 16'b1110110000010000;
            14'h5234: o_data_a = 16'b0000000000001110;
            14'h5235: o_data_a = 16'b1110001100001000;
            14'h5236: o_data_a = 16'b0101001000111010;
            14'h5237: o_data_a = 16'b1110110000010000;
            14'h5238: o_data_a = 16'b0000000001011111;
            14'h5239: o_data_a = 16'b1110101010000111;
            14'h523a: o_data_a = 16'b0000000000000000;
            14'h523b: o_data_a = 16'b1111110010101000;
            14'h523c: o_data_a = 16'b1111110000010000;
            14'h523d: o_data_a = 16'b0000000000000001;
            14'h523e: o_data_a = 16'b1111110000100000;
            14'h523f: o_data_a = 16'b1110001100001000;
            14'h5240: o_data_a = 16'b0000000000000010;
            14'h5241: o_data_a = 16'b1111110000100000;
            14'h5242: o_data_a = 16'b1111110000010000;
            14'h5243: o_data_a = 16'b0000000000000000;
            14'h5244: o_data_a = 16'b1111110111101000;
            14'h5245: o_data_a = 16'b1110110010100000;
            14'h5246: o_data_a = 16'b1110001100001000;
            14'h5247: o_data_a = 16'b0000000000000001;
            14'h5248: o_data_a = 16'b1111110000100000;
            14'h5249: o_data_a = 16'b1111110000010000;
            14'h524a: o_data_a = 16'b0000000000000000;
            14'h524b: o_data_a = 16'b1111110111101000;
            14'h524c: o_data_a = 16'b1110110010100000;
            14'h524d: o_data_a = 16'b1110001100001000;
            14'h524e: o_data_a = 16'b0000000000010000;
            14'h524f: o_data_a = 16'b1110110000010000;
            14'h5250: o_data_a = 16'b0000000000000000;
            14'h5251: o_data_a = 16'b1111110111101000;
            14'h5252: o_data_a = 16'b1110110010100000;
            14'h5253: o_data_a = 16'b1110001100001000;
            14'h5254: o_data_a = 16'b0000000000000010;
            14'h5255: o_data_a = 16'b1110110000010000;
            14'h5256: o_data_a = 16'b0000000000001101;
            14'h5257: o_data_a = 16'b1110001100001000;
            14'h5258: o_data_a = 16'b0001101010100110;
            14'h5259: o_data_a = 16'b1110110000010000;
            14'h525a: o_data_a = 16'b0000000000001110;
            14'h525b: o_data_a = 16'b1110001100001000;
            14'h525c: o_data_a = 16'b0101001001100000;
            14'h525d: o_data_a = 16'b1110110000010000;
            14'h525e: o_data_a = 16'b0000000001011111;
            14'h525f: o_data_a = 16'b1110101010000111;
            14'h5260: o_data_a = 16'b0000000000000000;
            14'h5261: o_data_a = 16'b1111110010101000;
            14'h5262: o_data_a = 16'b1111110000010000;
            14'h5263: o_data_a = 16'b1110110010100000;
            14'h5264: o_data_a = 16'b1111000111001000;
            14'h5265: o_data_a = 16'b0000000000000000;
            14'h5266: o_data_a = 16'b1111110010101000;
            14'h5267: o_data_a = 16'b1111110000010000;
            14'h5268: o_data_a = 16'b0000000000000001;
            14'h5269: o_data_a = 16'b1111110111100000;
            14'h526a: o_data_a = 16'b1110001100001000;
            14'h526b: o_data_a = 16'b0000000000000010;
            14'h526c: o_data_a = 16'b1111110111100000;
            14'h526d: o_data_a = 16'b1111110000010000;
            14'h526e: o_data_a = 16'b0000000000000000;
            14'h526f: o_data_a = 16'b1111110111101000;
            14'h5270: o_data_a = 16'b1110110010100000;
            14'h5271: o_data_a = 16'b1110001100001000;
            14'h5272: o_data_a = 16'b0000000000100000;
            14'h5273: o_data_a = 16'b1110110000010000;
            14'h5274: o_data_a = 16'b0000000000000000;
            14'h5275: o_data_a = 16'b1111110111101000;
            14'h5276: o_data_a = 16'b1110110010100000;
            14'h5277: o_data_a = 16'b1110001100001000;
            14'h5278: o_data_a = 16'b0000000000000010;
            14'h5279: o_data_a = 16'b1110110000010000;
            14'h527a: o_data_a = 16'b0000000000001101;
            14'h527b: o_data_a = 16'b1110001100001000;
            14'h527c: o_data_a = 16'b0001101010100110;
            14'h527d: o_data_a = 16'b1110110000010000;
            14'h527e: o_data_a = 16'b0000000000001110;
            14'h527f: o_data_a = 16'b1110001100001000;
            14'h5280: o_data_a = 16'b0101001010000100;
            14'h5281: o_data_a = 16'b1110110000010000;
            14'h5282: o_data_a = 16'b0000000001011111;
            14'h5283: o_data_a = 16'b1110101010000111;
            14'h5284: o_data_a = 16'b0000000000000001;
            14'h5285: o_data_a = 16'b1111110000100000;
            14'h5286: o_data_a = 16'b1111110000010000;
            14'h5287: o_data_a = 16'b0000000000000000;
            14'h5288: o_data_a = 16'b1111110111101000;
            14'h5289: o_data_a = 16'b1110110010100000;
            14'h528a: o_data_a = 16'b1110001100001000;
            14'h528b: o_data_a = 16'b0000000000000000;
            14'h528c: o_data_a = 16'b1111110010101000;
            14'h528d: o_data_a = 16'b1111110000010000;
            14'h528e: o_data_a = 16'b1110110010100000;
            14'h528f: o_data_a = 16'b1111000010001000;
            14'h5290: o_data_a = 16'b0000000000000000;
            14'h5291: o_data_a = 16'b1111110010101000;
            14'h5292: o_data_a = 16'b1111110000010000;
            14'h5293: o_data_a = 16'b0000000000000001;
            14'h5294: o_data_a = 16'b1111110111100000;
            14'h5295: o_data_a = 16'b1110110111100000;
            14'h5296: o_data_a = 16'b1110001100001000;
            14'h5297: o_data_a = 16'b0000000000000001;
            14'h5298: o_data_a = 16'b1111110111100000;
            14'h5299: o_data_a = 16'b1110110111100000;
            14'h529a: o_data_a = 16'b1111110000010000;
            14'h529b: o_data_a = 16'b0000000000000000;
            14'h529c: o_data_a = 16'b1111110111101000;
            14'h529d: o_data_a = 16'b1110110010100000;
            14'h529e: o_data_a = 16'b1110001100001000;
            14'h529f: o_data_a = 16'b0000000000000001;
            14'h52a0: o_data_a = 16'b1111110111100000;
            14'h52a1: o_data_a = 16'b1111110000010000;
            14'h52a2: o_data_a = 16'b0000000000000000;
            14'h52a3: o_data_a = 16'b1111110111101000;
            14'h52a4: o_data_a = 16'b1110110010100000;
            14'h52a5: o_data_a = 16'b1110001100001000;
            14'h52a6: o_data_a = 16'b0000000000011101;
            14'h52a7: o_data_a = 16'b1111110000010000;
            14'h52a8: o_data_a = 16'b0000000000000000;
            14'h52a9: o_data_a = 16'b1111110111101000;
            14'h52aa: o_data_a = 16'b1110110010100000;
            14'h52ab: o_data_a = 16'b1110001100001000;
            14'h52ac: o_data_a = 16'b0000000000000000;
            14'h52ad: o_data_a = 16'b1111110010101000;
            14'h52ae: o_data_a = 16'b1111110000010000;
            14'h52af: o_data_a = 16'b1110110010100000;
            14'h52b0: o_data_a = 16'b1111000010001000;
            14'h52b1: o_data_a = 16'b0000000000000000;
            14'h52b2: o_data_a = 16'b1111110010101000;
            14'h52b3: o_data_a = 16'b1111110000010000;
            14'h52b4: o_data_a = 16'b0000000000000100;
            14'h52b5: o_data_a = 16'b1110001100001000;
            14'h52b6: o_data_a = 16'b0000000000000100;
            14'h52b7: o_data_a = 16'b1111110000100000;
            14'h52b8: o_data_a = 16'b1111110000010000;
            14'h52b9: o_data_a = 16'b0000000000000000;
            14'h52ba: o_data_a = 16'b1111110111101000;
            14'h52bb: o_data_a = 16'b1110110010100000;
            14'h52bc: o_data_a = 16'b1110001100001000;
            14'h52bd: o_data_a = 16'b0000000000000010;
            14'h52be: o_data_a = 16'b1110110000010000;
            14'h52bf: o_data_a = 16'b0000000000001101;
            14'h52c0: o_data_a = 16'b1110001100001000;
            14'h52c1: o_data_a = 16'b0101000011011101;
            14'h52c2: o_data_a = 16'b1110110000010000;
            14'h52c3: o_data_a = 16'b0000000000001110;
            14'h52c4: o_data_a = 16'b1110001100001000;
            14'h52c5: o_data_a = 16'b0101001011001001;
            14'h52c6: o_data_a = 16'b1110110000010000;
            14'h52c7: o_data_a = 16'b0000000001011111;
            14'h52c8: o_data_a = 16'b1110101010000111;
            14'h52c9: o_data_a = 16'b0000000000000000;
            14'h52ca: o_data_a = 16'b1111110010101000;
            14'h52cb: o_data_a = 16'b1111110000010000;
            14'h52cc: o_data_a = 16'b0000000000000101;
            14'h52cd: o_data_a = 16'b1110001100001000;
            14'h52ce: o_data_a = 16'b0000000000000000;
            14'h52cf: o_data_a = 16'b1111110111001000;
            14'h52d0: o_data_a = 16'b1111110010100000;
            14'h52d1: o_data_a = 16'b1110101010001000;
            14'h52d2: o_data_a = 16'b0000000000110110;
            14'h52d3: o_data_a = 16'b1110101010000111;
            14'h52d4: o_data_a = 16'b0000000000000010;
            14'h52d5: o_data_a = 16'b1111110111100000;
            14'h52d6: o_data_a = 16'b1110110111100000;
            14'h52d7: o_data_a = 16'b1111110000010000;
            14'h52d8: o_data_a = 16'b0000000000000000;
            14'h52d9: o_data_a = 16'b1111110111101000;
            14'h52da: o_data_a = 16'b1110110010100000;
            14'h52db: o_data_a = 16'b1110001100001000;
            14'h52dc: o_data_a = 16'b0000000000000000;
            14'h52dd: o_data_a = 16'b1111110010101000;
            14'h52de: o_data_a = 16'b1111110000010000;
            14'h52df: o_data_a = 16'b0101001011100011;
            14'h52e0: o_data_a = 16'b1110001100000101;
            14'h52e1: o_data_a = 16'b0101001100000100;
            14'h52e2: o_data_a = 16'b1110101010000111;
            14'h52e3: o_data_a = 16'b0000000000000010;
            14'h52e4: o_data_a = 16'b1111110111100000;
            14'h52e5: o_data_a = 16'b1111110000010000;
            14'h52e6: o_data_a = 16'b0000000000000000;
            14'h52e7: o_data_a = 16'b1111110111101000;
            14'h52e8: o_data_a = 16'b1110110010100000;
            14'h52e9: o_data_a = 16'b1110001100001000;
            14'h52ea: o_data_a = 16'b0000000000000010;
            14'h52eb: o_data_a = 16'b1111110000100000;
            14'h52ec: o_data_a = 16'b1111110000010000;
            14'h52ed: o_data_a = 16'b0000000000000000;
            14'h52ee: o_data_a = 16'b1111110111101000;
            14'h52ef: o_data_a = 16'b1110110010100000;
            14'h52f0: o_data_a = 16'b1110001100001000;
            14'h52f1: o_data_a = 16'b0000000000000010;
            14'h52f2: o_data_a = 16'b1110110000010000;
            14'h52f3: o_data_a = 16'b0000000000001101;
            14'h52f4: o_data_a = 16'b1110001100001000;
            14'h52f5: o_data_a = 16'b0101000110101011;
            14'h52f6: o_data_a = 16'b1110110000010000;
            14'h52f7: o_data_a = 16'b0000000000001110;
            14'h52f8: o_data_a = 16'b1110001100001000;
            14'h52f9: o_data_a = 16'b0101001011111101;
            14'h52fa: o_data_a = 16'b1110110000010000;
            14'h52fb: o_data_a = 16'b0000000001011111;
            14'h52fc: o_data_a = 16'b1110101010000111;
            14'h52fd: o_data_a = 16'b0000000000000000;
            14'h52fe: o_data_a = 16'b1111110010101000;
            14'h52ff: o_data_a = 16'b1111110000010000;
            14'h5300: o_data_a = 16'b0000000000000101;
            14'h5301: o_data_a = 16'b1110001100001000;
            14'h5302: o_data_a = 16'b0101001100100011;
            14'h5303: o_data_a = 16'b1110101010000111;
            14'h5304: o_data_a = 16'b0000000000000010;
            14'h5305: o_data_a = 16'b1111110000100000;
            14'h5306: o_data_a = 16'b1111110000010000;
            14'h5307: o_data_a = 16'b0000000000000000;
            14'h5308: o_data_a = 16'b1111110111101000;
            14'h5309: o_data_a = 16'b1110110010100000;
            14'h530a: o_data_a = 16'b1110001100001000;
            14'h530b: o_data_a = 16'b0000000000000010;
            14'h530c: o_data_a = 16'b1111110111100000;
            14'h530d: o_data_a = 16'b1111110000010000;
            14'h530e: o_data_a = 16'b0000000000000000;
            14'h530f: o_data_a = 16'b1111110111101000;
            14'h5310: o_data_a = 16'b1110110010100000;
            14'h5311: o_data_a = 16'b1110001100001000;
            14'h5312: o_data_a = 16'b0000000000000010;
            14'h5313: o_data_a = 16'b1110110000010000;
            14'h5314: o_data_a = 16'b0000000000001101;
            14'h5315: o_data_a = 16'b1110001100001000;
            14'h5316: o_data_a = 16'b0101000110101011;
            14'h5317: o_data_a = 16'b1110110000010000;
            14'h5318: o_data_a = 16'b0000000000001110;
            14'h5319: o_data_a = 16'b1110001100001000;
            14'h531a: o_data_a = 16'b0101001100011110;
            14'h531b: o_data_a = 16'b1110110000010000;
            14'h531c: o_data_a = 16'b0000000001011111;
            14'h531d: o_data_a = 16'b1110101010000111;
            14'h531e: o_data_a = 16'b0000000000000000;
            14'h531f: o_data_a = 16'b1111110010101000;
            14'h5320: o_data_a = 16'b1111110000010000;
            14'h5321: o_data_a = 16'b0000000000000101;
            14'h5322: o_data_a = 16'b1110001100001000;
            14'h5323: o_data_a = 16'b0000000000000000;
            14'h5324: o_data_a = 16'b1111110111001000;
            14'h5325: o_data_a = 16'b1111110010100000;
            14'h5326: o_data_a = 16'b1110101010001000;
            14'h5327: o_data_a = 16'b0000000000110110;
            14'h5328: o_data_a = 16'b1110101010000111;
            14'h5329: o_data_a = 16'b0000000000001011;
            14'h532a: o_data_a = 16'b1110110000010000;
            14'h532b: o_data_a = 16'b1110001110010000;
            14'h532c: o_data_a = 16'b0000000000000000;
            14'h532d: o_data_a = 16'b1111110111101000;
            14'h532e: o_data_a = 16'b1110110010100000;
            14'h532f: o_data_a = 16'b1110101010001000;
            14'h5330: o_data_a = 16'b0101001100101011;
            14'h5331: o_data_a = 16'b1110001100000001;
            14'h5332: o_data_a = 16'b0000000000000010;
            14'h5333: o_data_a = 16'b1111110000100000;
            14'h5334: o_data_a = 16'b1111110000010000;
            14'h5335: o_data_a = 16'b0000000000000000;
            14'h5336: o_data_a = 16'b1111110111101000;
            14'h5337: o_data_a = 16'b1110110010100000;
            14'h5338: o_data_a = 16'b1110001100001000;
            14'h5339: o_data_a = 16'b0000000000000000;
            14'h533a: o_data_a = 16'b1111110111001000;
            14'h533b: o_data_a = 16'b1111110010100000;
            14'h533c: o_data_a = 16'b1110101010001000;
            14'h533d: o_data_a = 16'b0101001101000001;
            14'h533e: o_data_a = 16'b1110110000010000;
            14'h533f: o_data_a = 16'b0000000000100110;
            14'h5340: o_data_a = 16'b1110101010000111;
            14'h5341: o_data_a = 16'b0000000000000010;
            14'h5342: o_data_a = 16'b1111110111100000;
            14'h5343: o_data_a = 16'b1110110111100000;
            14'h5344: o_data_a = 16'b1111110000010000;
            14'h5345: o_data_a = 16'b0000000000000000;
            14'h5346: o_data_a = 16'b1111110111101000;
            14'h5347: o_data_a = 16'b1110110010100000;
            14'h5348: o_data_a = 16'b1110001100001000;
            14'h5349: o_data_a = 16'b0000000111111111;
            14'h534a: o_data_a = 16'b1110110000010000;
            14'h534b: o_data_a = 16'b0000000000000000;
            14'h534c: o_data_a = 16'b1111110111101000;
            14'h534d: o_data_a = 16'b1110110010100000;
            14'h534e: o_data_a = 16'b1110001100001000;
            14'h534f: o_data_a = 16'b0101001101010011;
            14'h5350: o_data_a = 16'b1110110000010000;
            14'h5351: o_data_a = 16'b0000000000010110;
            14'h5352: o_data_a = 16'b1110101010000111;
            14'h5353: o_data_a = 16'b0000000000000000;
            14'h5354: o_data_a = 16'b1111110010101000;
            14'h5355: o_data_a = 16'b1111110000010000;
            14'h5356: o_data_a = 16'b1110110010100000;
            14'h5357: o_data_a = 16'b1111010101001000;
            14'h5358: o_data_a = 16'b0000000000000010;
            14'h5359: o_data_a = 16'b1111110111100000;
            14'h535a: o_data_a = 16'b1111110000010000;
            14'h535b: o_data_a = 16'b0000000000000000;
            14'h535c: o_data_a = 16'b1111110111101000;
            14'h535d: o_data_a = 16'b1110110010100000;
            14'h535e: o_data_a = 16'b1110001100001000;
            14'h535f: o_data_a = 16'b0000000000000000;
            14'h5360: o_data_a = 16'b1111110111001000;
            14'h5361: o_data_a = 16'b1111110010100000;
            14'h5362: o_data_a = 16'b1110101010001000;
            14'h5363: o_data_a = 16'b0101001101100111;
            14'h5364: o_data_a = 16'b1110110000010000;
            14'h5365: o_data_a = 16'b0000000000100110;
            14'h5366: o_data_a = 16'b1110101010000111;
            14'h5367: o_data_a = 16'b0000000000000000;
            14'h5368: o_data_a = 16'b1111110010101000;
            14'h5369: o_data_a = 16'b1111110000010000;
            14'h536a: o_data_a = 16'b1110110010100000;
            14'h536b: o_data_a = 16'b1111010101001000;
            14'h536c: o_data_a = 16'b0000000000000010;
            14'h536d: o_data_a = 16'b1111110000010000;
            14'h536e: o_data_a = 16'b0000000000000011;
            14'h536f: o_data_a = 16'b1110000010100000;
            14'h5370: o_data_a = 16'b1111110000010000;
            14'h5371: o_data_a = 16'b0000000000000000;
            14'h5372: o_data_a = 16'b1111110111101000;
            14'h5373: o_data_a = 16'b1110110010100000;
            14'h5374: o_data_a = 16'b1110001100001000;
            14'h5375: o_data_a = 16'b0000000011111111;
            14'h5376: o_data_a = 16'b1110110000010000;
            14'h5377: o_data_a = 16'b0000000000000000;
            14'h5378: o_data_a = 16'b1111110111101000;
            14'h5379: o_data_a = 16'b1110110010100000;
            14'h537a: o_data_a = 16'b1110001100001000;
            14'h537b: o_data_a = 16'b0101001101111111;
            14'h537c: o_data_a = 16'b1110110000010000;
            14'h537d: o_data_a = 16'b0000000000010110;
            14'h537e: o_data_a = 16'b1110101010000111;
            14'h537f: o_data_a = 16'b0000000000000000;
            14'h5380: o_data_a = 16'b1111110010101000;
            14'h5381: o_data_a = 16'b1111110000010000;
            14'h5382: o_data_a = 16'b1110110010100000;
            14'h5383: o_data_a = 16'b1111010101001000;
            14'h5384: o_data_a = 16'b0000000000000000;
            14'h5385: o_data_a = 16'b1111110010101000;
            14'h5386: o_data_a = 16'b1111110000010000;
            14'h5387: o_data_a = 16'b0101001110001011;
            14'h5388: o_data_a = 16'b1110001100000101;
            14'h5389: o_data_a = 16'b0101001110100010;
            14'h538a: o_data_a = 16'b1110101010000111;
            14'h538b: o_data_a = 16'b0000000000001000;
            14'h538c: o_data_a = 16'b1110110000010000;
            14'h538d: o_data_a = 16'b0000000000000000;
            14'h538e: o_data_a = 16'b1111110111101000;
            14'h538f: o_data_a = 16'b1110110010100000;
            14'h5390: o_data_a = 16'b1110001100001000;
            14'h5391: o_data_a = 16'b0000000000000001;
            14'h5392: o_data_a = 16'b1110110000010000;
            14'h5393: o_data_a = 16'b0000000000001101;
            14'h5394: o_data_a = 16'b1110001100001000;
            14'h5395: o_data_a = 16'b0110101011011001;
            14'h5396: o_data_a = 16'b1110110000010000;
            14'h5397: o_data_a = 16'b0000000000001110;
            14'h5398: o_data_a = 16'b1110001100001000;
            14'h5399: o_data_a = 16'b0101001110011101;
            14'h539a: o_data_a = 16'b1110110000010000;
            14'h539b: o_data_a = 16'b0000000001011111;
            14'h539c: o_data_a = 16'b1110101010000111;
            14'h539d: o_data_a = 16'b0000000000000000;
            14'h539e: o_data_a = 16'b1111110010101000;
            14'h539f: o_data_a = 16'b1111110000010000;
            14'h53a0: o_data_a = 16'b0000000000000101;
            14'h53a1: o_data_a = 16'b1110001100001000;
            14'h53a2: o_data_a = 16'b0000000000000010;
            14'h53a3: o_data_a = 16'b1111110111100000;
            14'h53a4: o_data_a = 16'b1110110111100000;
            14'h53a5: o_data_a = 16'b1111110000010000;
            14'h53a6: o_data_a = 16'b0000000000000000;
            14'h53a7: o_data_a = 16'b1111110111101000;
            14'h53a8: o_data_a = 16'b1110110010100000;
            14'h53a9: o_data_a = 16'b1110001100001000;
            14'h53aa: o_data_a = 16'b0000000000000010;
            14'h53ab: o_data_a = 16'b1111110000100000;
            14'h53ac: o_data_a = 16'b1111110000010000;
            14'h53ad: o_data_a = 16'b0000000000000000;
            14'h53ae: o_data_a = 16'b1111110111101000;
            14'h53af: o_data_a = 16'b1110110010100000;
            14'h53b0: o_data_a = 16'b1110001100001000;
            14'h53b1: o_data_a = 16'b0000000000000000;
            14'h53b2: o_data_a = 16'b1111110010101000;
            14'h53b3: o_data_a = 16'b1111110000010000;
            14'h53b4: o_data_a = 16'b1110110010100000;
            14'h53b5: o_data_a = 16'b1111000111001000;
            14'h53b6: o_data_a = 16'b0000000000000001;
            14'h53b7: o_data_a = 16'b1110110000010000;
            14'h53b8: o_data_a = 16'b0000000000001101;
            14'h53b9: o_data_a = 16'b1110001100001000;
            14'h53ba: o_data_a = 16'b0001101001110110;
            14'h53bb: o_data_a = 16'b1110110000010000;
            14'h53bc: o_data_a = 16'b0000000000001110;
            14'h53bd: o_data_a = 16'b1110001100001000;
            14'h53be: o_data_a = 16'b0101001111000010;
            14'h53bf: o_data_a = 16'b1110110000010000;
            14'h53c0: o_data_a = 16'b0000000001011111;
            14'h53c1: o_data_a = 16'b1110101010000111;
            14'h53c2: o_data_a = 16'b0000000000000000;
            14'h53c3: o_data_a = 16'b1111110010101000;
            14'h53c4: o_data_a = 16'b1111110000010000;
            14'h53c5: o_data_a = 16'b0000000000000001;
            14'h53c6: o_data_a = 16'b1111110111100000;
            14'h53c7: o_data_a = 16'b1110110111100000;
            14'h53c8: o_data_a = 16'b1110110111100000;
            14'h53c9: o_data_a = 16'b1110001100001000;
            14'h53ca: o_data_a = 16'b0000000000000010;
            14'h53cb: o_data_a = 16'b1111110000010000;
            14'h53cc: o_data_a = 16'b0000000000000011;
            14'h53cd: o_data_a = 16'b1110000010100000;
            14'h53ce: o_data_a = 16'b1111110000010000;
            14'h53cf: o_data_a = 16'b0000000000000000;
            14'h53d0: o_data_a = 16'b1111110111101000;
            14'h53d1: o_data_a = 16'b1110110010100000;
            14'h53d2: o_data_a = 16'b1110001100001000;
            14'h53d3: o_data_a = 16'b0000000000000010;
            14'h53d4: o_data_a = 16'b1111110111100000;
            14'h53d5: o_data_a = 16'b1111110000010000;
            14'h53d6: o_data_a = 16'b0000000000000000;
            14'h53d7: o_data_a = 16'b1111110111101000;
            14'h53d8: o_data_a = 16'b1110110010100000;
            14'h53d9: o_data_a = 16'b1110001100001000;
            14'h53da: o_data_a = 16'b0000000000000000;
            14'h53db: o_data_a = 16'b1111110010101000;
            14'h53dc: o_data_a = 16'b1111110000010000;
            14'h53dd: o_data_a = 16'b1110110010100000;
            14'h53de: o_data_a = 16'b1111000111001000;
            14'h53df: o_data_a = 16'b0000000000000001;
            14'h53e0: o_data_a = 16'b1110110000010000;
            14'h53e1: o_data_a = 16'b0000000000001101;
            14'h53e2: o_data_a = 16'b1110001100001000;
            14'h53e3: o_data_a = 16'b0001101001110110;
            14'h53e4: o_data_a = 16'b1110110000010000;
            14'h53e5: o_data_a = 16'b0000000000001110;
            14'h53e6: o_data_a = 16'b1110001100001000;
            14'h53e7: o_data_a = 16'b0101001111101011;
            14'h53e8: o_data_a = 16'b1110110000010000;
            14'h53e9: o_data_a = 16'b0000000001011111;
            14'h53ea: o_data_a = 16'b1110101010000111;
            14'h53eb: o_data_a = 16'b0000000000000000;
            14'h53ec: o_data_a = 16'b1111110010101000;
            14'h53ed: o_data_a = 16'b1111110000010000;
            14'h53ee: o_data_a = 16'b0000000000000001;
            14'h53ef: o_data_a = 16'b1111110111100000;
            14'h53f0: o_data_a = 16'b1110110111100000;
            14'h53f1: o_data_a = 16'b1110001100001000;
            14'h53f2: o_data_a = 16'b0000000000000001;
            14'h53f3: o_data_a = 16'b1111110000010000;
            14'h53f4: o_data_a = 16'b0000000000000011;
            14'h53f5: o_data_a = 16'b1110000010100000;
            14'h53f6: o_data_a = 16'b1111110000010000;
            14'h53f7: o_data_a = 16'b0000000000000000;
            14'h53f8: o_data_a = 16'b1111110111101000;
            14'h53f9: o_data_a = 16'b1110110010100000;
            14'h53fa: o_data_a = 16'b1110001100001000;
            14'h53fb: o_data_a = 16'b0000000000000001;
            14'h53fc: o_data_a = 16'b1111110111100000;
            14'h53fd: o_data_a = 16'b1110110111100000;
            14'h53fe: o_data_a = 16'b1111110000010000;
            14'h53ff: o_data_a = 16'b0000000000000000;
            14'h5400: o_data_a = 16'b1111110111101000;
            14'h5401: o_data_a = 16'b1110110010100000;
            14'h5402: o_data_a = 16'b1110001100001000;
            14'h5403: o_data_a = 16'b0101010000000111;
            14'h5404: o_data_a = 16'b1110110000010000;
            14'h5405: o_data_a = 16'b0000000000100110;
            14'h5406: o_data_a = 16'b1110101010000111;
            14'h5407: o_data_a = 16'b0000000000000000;
            14'h5408: o_data_a = 16'b1111110010101000;
            14'h5409: o_data_a = 16'b1111110000010000;
            14'h540a: o_data_a = 16'b0000000000000001;
            14'h540b: o_data_a = 16'b1111110111100000;
            14'h540c: o_data_a = 16'b1110110111100000;
            14'h540d: o_data_a = 16'b1110110111100000;
            14'h540e: o_data_a = 16'b1110110111100000;
            14'h540f: o_data_a = 16'b1110110111100000;
            14'h5410: o_data_a = 16'b1110110111100000;
            14'h5411: o_data_a = 16'b1110001100001000;
            14'h5412: o_data_a = 16'b0000000000000001;
            14'h5413: o_data_a = 16'b1111110000010000;
            14'h5414: o_data_a = 16'b0000000000000110;
            14'h5415: o_data_a = 16'b1110000010100000;
            14'h5416: o_data_a = 16'b1111110000010000;
            14'h5417: o_data_a = 16'b0000000000000000;
            14'h5418: o_data_a = 16'b1111110111101000;
            14'h5419: o_data_a = 16'b1110110010100000;
            14'h541a: o_data_a = 16'b1110001100001000;
            14'h541b: o_data_a = 16'b0000000000000010;
            14'h541c: o_data_a = 16'b1111110000010000;
            14'h541d: o_data_a = 16'b0000000000000011;
            14'h541e: o_data_a = 16'b1110000010100000;
            14'h541f: o_data_a = 16'b1111110000010000;
            14'h5420: o_data_a = 16'b0000000000000000;
            14'h5421: o_data_a = 16'b1111110111101000;
            14'h5422: o_data_a = 16'b1110110010100000;
            14'h5423: o_data_a = 16'b1110001100001000;
            14'h5424: o_data_a = 16'b0000000000000010;
            14'h5425: o_data_a = 16'b1111110111100000;
            14'h5426: o_data_a = 16'b1111110000010000;
            14'h5427: o_data_a = 16'b0000000000000000;
            14'h5428: o_data_a = 16'b1111110111101000;
            14'h5429: o_data_a = 16'b1110110010100000;
            14'h542a: o_data_a = 16'b1110001100001000;
            14'h542b: o_data_a = 16'b0101010000101111;
            14'h542c: o_data_a = 16'b1110110000010000;
            14'h542d: o_data_a = 16'b0000000000100110;
            14'h542e: o_data_a = 16'b1110101010000111;
            14'h542f: o_data_a = 16'b0000000000000000;
            14'h5430: o_data_a = 16'b1111110010101000;
            14'h5431: o_data_a = 16'b1111110000010000;
            14'h5432: o_data_a = 16'b1110110010100000;
            14'h5433: o_data_a = 16'b1111000000001000;
            14'h5434: o_data_a = 16'b0000000000000001;
            14'h5435: o_data_a = 16'b1111110000010000;
            14'h5436: o_data_a = 16'b0000000000000110;
            14'h5437: o_data_a = 16'b1110000010100000;
            14'h5438: o_data_a = 16'b1111110000010000;
            14'h5439: o_data_a = 16'b0000000000000000;
            14'h543a: o_data_a = 16'b1111110111101000;
            14'h543b: o_data_a = 16'b1110110010100000;
            14'h543c: o_data_a = 16'b1110001100001000;
            14'h543d: o_data_a = 16'b0000000000000000;
            14'h543e: o_data_a = 16'b1111110010100000;
            14'h543f: o_data_a = 16'b1111110001001000;
            14'h5440: o_data_a = 16'b0000000000000010;
            14'h5441: o_data_a = 16'b1111110111100000;
            14'h5442: o_data_a = 16'b1110110111100000;
            14'h5443: o_data_a = 16'b1111110000010000;
            14'h5444: o_data_a = 16'b0000000000000000;
            14'h5445: o_data_a = 16'b1111110111101000;
            14'h5446: o_data_a = 16'b1110110010100000;
            14'h5447: o_data_a = 16'b1110001100001000;
            14'h5448: o_data_a = 16'b0000000000000010;
            14'h5449: o_data_a = 16'b1111110000100000;
            14'h544a: o_data_a = 16'b1111110000010000;
            14'h544b: o_data_a = 16'b0000000000000000;
            14'h544c: o_data_a = 16'b1111110111101000;
            14'h544d: o_data_a = 16'b1110110010100000;
            14'h544e: o_data_a = 16'b1110001100001000;
            14'h544f: o_data_a = 16'b0101010001010011;
            14'h5450: o_data_a = 16'b1110110000010000;
            14'h5451: o_data_a = 16'b0000000000100110;
            14'h5452: o_data_a = 16'b1110101010000111;
            14'h5453: o_data_a = 16'b0000000000000000;
            14'h5454: o_data_a = 16'b1111110010101000;
            14'h5455: o_data_a = 16'b1111110000010000;
            14'h5456: o_data_a = 16'b1110110010100000;
            14'h5457: o_data_a = 16'b1111000000001000;
            14'h5458: o_data_a = 16'b0000000000000000;
            14'h5459: o_data_a = 16'b1111110010101000;
            14'h545a: o_data_a = 16'b1111110000010000;
            14'h545b: o_data_a = 16'b1110110010100000;
            14'h545c: o_data_a = 16'b1111010101001000;
            14'h545d: o_data_a = 16'b0000000000000000;
            14'h545e: o_data_a = 16'b1111110010101000;
            14'h545f: o_data_a = 16'b1111110000010000;
            14'h5460: o_data_a = 16'b0101010001100100;
            14'h5461: o_data_a = 16'b1110001100000101;
            14'h5462: o_data_a = 16'b0101010011000010;
            14'h5463: o_data_a = 16'b1110101010000111;
            14'h5464: o_data_a = 16'b0000000000000010;
            14'h5465: o_data_a = 16'b1111110000100000;
            14'h5466: o_data_a = 16'b1111110000010000;
            14'h5467: o_data_a = 16'b0000000000000000;
            14'h5468: o_data_a = 16'b1111110111101000;
            14'h5469: o_data_a = 16'b1110110010100000;
            14'h546a: o_data_a = 16'b1110001100001000;
            14'h546b: o_data_a = 16'b0000000000000000;
            14'h546c: o_data_a = 16'b1111110010101000;
            14'h546d: o_data_a = 16'b1111110000010000;
            14'h546e: o_data_a = 16'b0000000000000001;
            14'h546f: o_data_a = 16'b1111110111100000;
            14'h5470: o_data_a = 16'b1110110111100000;
            14'h5471: o_data_a = 16'b1110110111100000;
            14'h5472: o_data_a = 16'b1110110111100000;
            14'h5473: o_data_a = 16'b1110001100001000;
            14'h5474: o_data_a = 16'b0000000000000010;
            14'h5475: o_data_a = 16'b1111110111100000;
            14'h5476: o_data_a = 16'b1110110111100000;
            14'h5477: o_data_a = 16'b1111110000010000;
            14'h5478: o_data_a = 16'b0000000000000000;
            14'h5479: o_data_a = 16'b1111110111101000;
            14'h547a: o_data_a = 16'b1110110010100000;
            14'h547b: o_data_a = 16'b1110001100001000;
            14'h547c: o_data_a = 16'b0000000000000000;
            14'h547d: o_data_a = 16'b1111110010101000;
            14'h547e: o_data_a = 16'b1111110000010000;
            14'h547f: o_data_a = 16'b0000000000000010;
            14'h5480: o_data_a = 16'b1111110000100000;
            14'h5481: o_data_a = 16'b1110001100001000;
            14'h5482: o_data_a = 16'b0000000000000001;
            14'h5483: o_data_a = 16'b1111110000010000;
            14'h5484: o_data_a = 16'b0000000000000100;
            14'h5485: o_data_a = 16'b1110000010100000;
            14'h5486: o_data_a = 16'b1111110000010000;
            14'h5487: o_data_a = 16'b0000000000000000;
            14'h5488: o_data_a = 16'b1111110111101000;
            14'h5489: o_data_a = 16'b1110110010100000;
            14'h548a: o_data_a = 16'b1110001100001000;
            14'h548b: o_data_a = 16'b0000000000000000;
            14'h548c: o_data_a = 16'b1111110010101000;
            14'h548d: o_data_a = 16'b1111110000010000;
            14'h548e: o_data_a = 16'b0000000000000010;
            14'h548f: o_data_a = 16'b1111110111100000;
            14'h5490: o_data_a = 16'b1110110111100000;
            14'h5491: o_data_a = 16'b1110001100001000;
            14'h5492: o_data_a = 16'b0000000000000010;
            14'h5493: o_data_a = 16'b1111110111100000;
            14'h5494: o_data_a = 16'b1111110000010000;
            14'h5495: o_data_a = 16'b0000000000000000;
            14'h5496: o_data_a = 16'b1111110111101000;
            14'h5497: o_data_a = 16'b1110110010100000;
            14'h5498: o_data_a = 16'b1110001100001000;
            14'h5499: o_data_a = 16'b0000000000000000;
            14'h549a: o_data_a = 16'b1111110010101000;
            14'h549b: o_data_a = 16'b1111110000010000;
            14'h549c: o_data_a = 16'b0000000000000001;
            14'h549d: o_data_a = 16'b1111110111100000;
            14'h549e: o_data_a = 16'b1110110111100000;
            14'h549f: o_data_a = 16'b1110110111100000;
            14'h54a0: o_data_a = 16'b1110110111100000;
            14'h54a1: o_data_a = 16'b1110001100001000;
            14'h54a2: o_data_a = 16'b0000000000000010;
            14'h54a3: o_data_a = 16'b1111110000010000;
            14'h54a4: o_data_a = 16'b0000000000000011;
            14'h54a5: o_data_a = 16'b1110000010100000;
            14'h54a6: o_data_a = 16'b1111110000010000;
            14'h54a7: o_data_a = 16'b0000000000000000;
            14'h54a8: o_data_a = 16'b1111110111101000;
            14'h54a9: o_data_a = 16'b1110110010100000;
            14'h54aa: o_data_a = 16'b1110001100001000;
            14'h54ab: o_data_a = 16'b0000000000000000;
            14'h54ac: o_data_a = 16'b1111110010101000;
            14'h54ad: o_data_a = 16'b1111110000010000;
            14'h54ae: o_data_a = 16'b0000000000000010;
            14'h54af: o_data_a = 16'b1111110111100000;
            14'h54b0: o_data_a = 16'b1110001100001000;
            14'h54b1: o_data_a = 16'b0000000000000001;
            14'h54b2: o_data_a = 16'b1111110000010000;
            14'h54b3: o_data_a = 16'b0000000000000100;
            14'h54b4: o_data_a = 16'b1110000010100000;
            14'h54b5: o_data_a = 16'b1111110000010000;
            14'h54b6: o_data_a = 16'b0000000000000000;
            14'h54b7: o_data_a = 16'b1111110111101000;
            14'h54b8: o_data_a = 16'b1110110010100000;
            14'h54b9: o_data_a = 16'b1110001100001000;
            14'h54ba: o_data_a = 16'b0000000000000000;
            14'h54bb: o_data_a = 16'b1111110010101000;
            14'h54bc: o_data_a = 16'b1111110000010000;
            14'h54bd: o_data_a = 16'b0000000000000010;
            14'h54be: o_data_a = 16'b1111110111100000;
            14'h54bf: o_data_a = 16'b1110110111100000;
            14'h54c0: o_data_a = 16'b1110110111100000;
            14'h54c1: o_data_a = 16'b1110001100001000;
            14'h54c2: o_data_a = 16'b0000000000000001;
            14'h54c3: o_data_a = 16'b1111110000010000;
            14'h54c4: o_data_a = 16'b0000000000000110;
            14'h54c5: o_data_a = 16'b1110000010100000;
            14'h54c6: o_data_a = 16'b1111110000010000;
            14'h54c7: o_data_a = 16'b0000000000000000;
            14'h54c8: o_data_a = 16'b1111110111101000;
            14'h54c9: o_data_a = 16'b1110110010100000;
            14'h54ca: o_data_a = 16'b1110001100001000;
            14'h54cb: o_data_a = 16'b0000000000000000;
            14'h54cc: o_data_a = 16'b1111110010101000;
            14'h54cd: o_data_a = 16'b1111110000010000;
            14'h54ce: o_data_a = 16'b0101010011010010;
            14'h54cf: o_data_a = 16'b1110001100000101;
            14'h54d0: o_data_a = 16'b0101010101010100;
            14'h54d1: o_data_a = 16'b1110101010000111;
            14'h54d2: o_data_a = 16'b0000000000000001;
            14'h54d3: o_data_a = 16'b1111110000010000;
            14'h54d4: o_data_a = 16'b0000000000000011;
            14'h54d5: o_data_a = 16'b1110000010100000;
            14'h54d6: o_data_a = 16'b1111110000010000;
            14'h54d7: o_data_a = 16'b0000000000000000;
            14'h54d8: o_data_a = 16'b1111110111101000;
            14'h54d9: o_data_a = 16'b1110110010100000;
            14'h54da: o_data_a = 16'b1110001100001000;
            14'h54db: o_data_a = 16'b0000000000000000;
            14'h54dc: o_data_a = 16'b1111110010101000;
            14'h54dd: o_data_a = 16'b1111110000010000;
            14'h54de: o_data_a = 16'b0000000000000001;
            14'h54df: o_data_a = 16'b1111110111100000;
            14'h54e0: o_data_a = 16'b1110110111100000;
            14'h54e1: o_data_a = 16'b1110110111100000;
            14'h54e2: o_data_a = 16'b1110110111100000;
            14'h54e3: o_data_a = 16'b1110001100001000;
            14'h54e4: o_data_a = 16'b0000000000000001;
            14'h54e5: o_data_a = 16'b1111110111100000;
            14'h54e6: o_data_a = 16'b1110110111100000;
            14'h54e7: o_data_a = 16'b1111110000010000;
            14'h54e8: o_data_a = 16'b0000000000000000;
            14'h54e9: o_data_a = 16'b1111110111101000;
            14'h54ea: o_data_a = 16'b1110110010100000;
            14'h54eb: o_data_a = 16'b1110001100001000;
            14'h54ec: o_data_a = 16'b0000000000000000;
            14'h54ed: o_data_a = 16'b1111110010101000;
            14'h54ee: o_data_a = 16'b1111110000010000;
            14'h54ef: o_data_a = 16'b0000000000000001;
            14'h54f0: o_data_a = 16'b1111110111100000;
            14'h54f1: o_data_a = 16'b1110110111100000;
            14'h54f2: o_data_a = 16'b1110110111100000;
            14'h54f3: o_data_a = 16'b1110001100001000;
            14'h54f4: o_data_a = 16'b0000000000000001;
            14'h54f5: o_data_a = 16'b1111110000010000;
            14'h54f6: o_data_a = 16'b0000000000000100;
            14'h54f7: o_data_a = 16'b1110000010100000;
            14'h54f8: o_data_a = 16'b1111110000010000;
            14'h54f9: o_data_a = 16'b0000000000000000;
            14'h54fa: o_data_a = 16'b1111110111101000;
            14'h54fb: o_data_a = 16'b1110110010100000;
            14'h54fc: o_data_a = 16'b1110001100001000;
            14'h54fd: o_data_a = 16'b0000000000000000;
            14'h54fe: o_data_a = 16'b1111110010101000;
            14'h54ff: o_data_a = 16'b1111110000010000;
            14'h5500: o_data_a = 16'b0000000000000001;
            14'h5501: o_data_a = 16'b1111110111100000;
            14'h5502: o_data_a = 16'b1110110111100000;
            14'h5503: o_data_a = 16'b1110001100001000;
            14'h5504: o_data_a = 16'b0000000000000010;
            14'h5505: o_data_a = 16'b1111110111100000;
            14'h5506: o_data_a = 16'b1111110000010000;
            14'h5507: o_data_a = 16'b0000000000000000;
            14'h5508: o_data_a = 16'b1111110111101000;
            14'h5509: o_data_a = 16'b1110110010100000;
            14'h550a: o_data_a = 16'b1110001100001000;
            14'h550b: o_data_a = 16'b0000000000000000;
            14'h550c: o_data_a = 16'b1111110010101000;
            14'h550d: o_data_a = 16'b1111110000010000;
            14'h550e: o_data_a = 16'b0000000000000001;
            14'h550f: o_data_a = 16'b1111110111100000;
            14'h5510: o_data_a = 16'b1110001100001000;
            14'h5511: o_data_a = 16'b0000000000000010;
            14'h5512: o_data_a = 16'b1111110000100000;
            14'h5513: o_data_a = 16'b1111110000010000;
            14'h5514: o_data_a = 16'b0000000000000000;
            14'h5515: o_data_a = 16'b1111110111101000;
            14'h5516: o_data_a = 16'b1110110010100000;
            14'h5517: o_data_a = 16'b1110001100001000;
            14'h5518: o_data_a = 16'b0000000000000000;
            14'h5519: o_data_a = 16'b1111110010101000;
            14'h551a: o_data_a = 16'b1111110000010000;
            14'h551b: o_data_a = 16'b0000000000000001;
            14'h551c: o_data_a = 16'b1111110000100000;
            14'h551d: o_data_a = 16'b1110001100001000;
            14'h551e: o_data_a = 16'b0000000000000010;
            14'h551f: o_data_a = 16'b1111110000010000;
            14'h5520: o_data_a = 16'b0000000000000011;
            14'h5521: o_data_a = 16'b1110000010100000;
            14'h5522: o_data_a = 16'b1111110000010000;
            14'h5523: o_data_a = 16'b0000000000000000;
            14'h5524: o_data_a = 16'b1111110111101000;
            14'h5525: o_data_a = 16'b1110110010100000;
            14'h5526: o_data_a = 16'b1110001100001000;
            14'h5527: o_data_a = 16'b0000000000000001;
            14'h5528: o_data_a = 16'b1111110000010000;
            14'h5529: o_data_a = 16'b0000000000001000;
            14'h552a: o_data_a = 16'b1110000010010000;
            14'h552b: o_data_a = 16'b0000000000001101;
            14'h552c: o_data_a = 16'b1110001100001000;
            14'h552d: o_data_a = 16'b0000000000000000;
            14'h552e: o_data_a = 16'b1111110010101000;
            14'h552f: o_data_a = 16'b1111110000010000;
            14'h5530: o_data_a = 16'b0000000000001101;
            14'h5531: o_data_a = 16'b1111110000100000;
            14'h5532: o_data_a = 16'b1110001100001000;
            14'h5533: o_data_a = 16'b0000000000000010;
            14'h5534: o_data_a = 16'b1111110000100000;
            14'h5535: o_data_a = 16'b1111110000010000;
            14'h5536: o_data_a = 16'b0000000000000000;
            14'h5537: o_data_a = 16'b1111110111101000;
            14'h5538: o_data_a = 16'b1110110010100000;
            14'h5539: o_data_a = 16'b1110001100001000;
            14'h553a: o_data_a = 16'b0000000000000010;
            14'h553b: o_data_a = 16'b1111110111100000;
            14'h553c: o_data_a = 16'b1110110111100000;
            14'h553d: o_data_a = 16'b1111110000010000;
            14'h553e: o_data_a = 16'b0000000000000000;
            14'h553f: o_data_a = 16'b1111110111101000;
            14'h5540: o_data_a = 16'b1110110010100000;
            14'h5541: o_data_a = 16'b1110001100001000;
            14'h5542: o_data_a = 16'b0101010101000110;
            14'h5543: o_data_a = 16'b1110110000010000;
            14'h5544: o_data_a = 16'b0000000000010110;
            14'h5545: o_data_a = 16'b1110101010000111;
            14'h5546: o_data_a = 16'b0000000000000001;
            14'h5547: o_data_a = 16'b1111110000010000;
            14'h5548: o_data_a = 16'b0000000000000111;
            14'h5549: o_data_a = 16'b1110000010010000;
            14'h554a: o_data_a = 16'b0000000000001101;
            14'h554b: o_data_a = 16'b1110001100001000;
            14'h554c: o_data_a = 16'b0000000000000000;
            14'h554d: o_data_a = 16'b1111110010101000;
            14'h554e: o_data_a = 16'b1111110000010000;
            14'h554f: o_data_a = 16'b0000000000001101;
            14'h5550: o_data_a = 16'b1111110000100000;
            14'h5551: o_data_a = 16'b1110001100001000;
            14'h5552: o_data_a = 16'b0101010110100010;
            14'h5553: o_data_a = 16'b1110101010000111;
            14'h5554: o_data_a = 16'b0000000000000010;
            14'h5555: o_data_a = 16'b1111110000100000;
            14'h5556: o_data_a = 16'b1111110000010000;
            14'h5557: o_data_a = 16'b0000000000000000;
            14'h5558: o_data_a = 16'b1111110111101000;
            14'h5559: o_data_a = 16'b1110110010100000;
            14'h555a: o_data_a = 16'b1110001100001000;
            14'h555b: o_data_a = 16'b0000000000000000;
            14'h555c: o_data_a = 16'b1111110010101000;
            14'h555d: o_data_a = 16'b1111110000010000;
            14'h555e: o_data_a = 16'b0000000000000001;
            14'h555f: o_data_a = 16'b1111110111100000;
            14'h5560: o_data_a = 16'b1110001100001000;
            14'h5561: o_data_a = 16'b0000000000000010;
            14'h5562: o_data_a = 16'b1111110111100000;
            14'h5563: o_data_a = 16'b1111110000010000;
            14'h5564: o_data_a = 16'b0000000000000000;
            14'h5565: o_data_a = 16'b1111110111101000;
            14'h5566: o_data_a = 16'b1110110010100000;
            14'h5567: o_data_a = 16'b1110001100001000;
            14'h5568: o_data_a = 16'b0000000000000000;
            14'h5569: o_data_a = 16'b1111110010101000;
            14'h556a: o_data_a = 16'b1111110000010000;
            14'h556b: o_data_a = 16'b0000000000000001;
            14'h556c: o_data_a = 16'b1111110000100000;
            14'h556d: o_data_a = 16'b1110001100001000;
            14'h556e: o_data_a = 16'b0000000000000010;
            14'h556f: o_data_a = 16'b1111110111100000;
            14'h5570: o_data_a = 16'b1110110111100000;
            14'h5571: o_data_a = 16'b1111110000010000;
            14'h5572: o_data_a = 16'b0000000000000000;
            14'h5573: o_data_a = 16'b1111110111101000;
            14'h5574: o_data_a = 16'b1110110010100000;
            14'h5575: o_data_a = 16'b1110001100001000;
            14'h5576: o_data_a = 16'b0000000000000001;
            14'h5577: o_data_a = 16'b1111110000010000;
            14'h5578: o_data_a = 16'b0000000000001000;
            14'h5579: o_data_a = 16'b1110000010010000;
            14'h557a: o_data_a = 16'b0000000000001101;
            14'h557b: o_data_a = 16'b1110001100001000;
            14'h557c: o_data_a = 16'b0000000000000000;
            14'h557d: o_data_a = 16'b1111110010101000;
            14'h557e: o_data_a = 16'b1111110000010000;
            14'h557f: o_data_a = 16'b0000000000001101;
            14'h5580: o_data_a = 16'b1111110000100000;
            14'h5581: o_data_a = 16'b1110001100001000;
            14'h5582: o_data_a = 16'b0000000000000010;
            14'h5583: o_data_a = 16'b1111110111100000;
            14'h5584: o_data_a = 16'b1111110000010000;
            14'h5585: o_data_a = 16'b0000000000000000;
            14'h5586: o_data_a = 16'b1111110111101000;
            14'h5587: o_data_a = 16'b1110110010100000;
            14'h5588: o_data_a = 16'b1110001100001000;
            14'h5589: o_data_a = 16'b0000000000000010;
            14'h558a: o_data_a = 16'b1111110000010000;
            14'h558b: o_data_a = 16'b0000000000000011;
            14'h558c: o_data_a = 16'b1110000010100000;
            14'h558d: o_data_a = 16'b1111110000010000;
            14'h558e: o_data_a = 16'b0000000000000000;
            14'h558f: o_data_a = 16'b1111110111101000;
            14'h5590: o_data_a = 16'b1110110010100000;
            14'h5591: o_data_a = 16'b1110001100001000;
            14'h5592: o_data_a = 16'b0101010110010110;
            14'h5593: o_data_a = 16'b1110110000010000;
            14'h5594: o_data_a = 16'b0000000000010110;
            14'h5595: o_data_a = 16'b1110101010000111;
            14'h5596: o_data_a = 16'b0000000000000001;
            14'h5597: o_data_a = 16'b1111110000010000;
            14'h5598: o_data_a = 16'b0000000000000111;
            14'h5599: o_data_a = 16'b1110000010010000;
            14'h559a: o_data_a = 16'b0000000000001101;
            14'h559b: o_data_a = 16'b1110001100001000;
            14'h559c: o_data_a = 16'b0000000000000000;
            14'h559d: o_data_a = 16'b1111110010101000;
            14'h559e: o_data_a = 16'b1111110000010000;
            14'h559f: o_data_a = 16'b0000000000001101;
            14'h55a0: o_data_a = 16'b1111110000100000;
            14'h55a1: o_data_a = 16'b1110001100001000;
            14'h55a2: o_data_a = 16'b0000000000000010;
            14'h55a3: o_data_a = 16'b1110110000010000;
            14'h55a4: o_data_a = 16'b0000000000000000;
            14'h55a5: o_data_a = 16'b1111110111101000;
            14'h55a6: o_data_a = 16'b1110110010100000;
            14'h55a7: o_data_a = 16'b1110001100001000;
            14'h55a8: o_data_a = 16'b0000000000000001;
            14'h55a9: o_data_a = 16'b1111110111100000;
            14'h55aa: o_data_a = 16'b1110110111100000;
            14'h55ab: o_data_a = 16'b1111110000010000;
            14'h55ac: o_data_a = 16'b0000000000000000;
            14'h55ad: o_data_a = 16'b1111110111101000;
            14'h55ae: o_data_a = 16'b1110110010100000;
            14'h55af: o_data_a = 16'b1110001100001000;
            14'h55b0: o_data_a = 16'b0000000000000010;
            14'h55b1: o_data_a = 16'b1110110000010000;
            14'h55b2: o_data_a = 16'b0000000000001101;
            14'h55b3: o_data_a = 16'b1110001100001000;
            14'h55b4: o_data_a = 16'b0001101010100110;
            14'h55b5: o_data_a = 16'b1110110000010000;
            14'h55b6: o_data_a = 16'b0000000000001110;
            14'h55b7: o_data_a = 16'b1110001100001000;
            14'h55b8: o_data_a = 16'b0101010110111100;
            14'h55b9: o_data_a = 16'b1110110000010000;
            14'h55ba: o_data_a = 16'b0000000001011111;
            14'h55bb: o_data_a = 16'b1110101010000111;
            14'h55bc: o_data_a = 16'b0000000000000001;
            14'h55bd: o_data_a = 16'b1111110000010000;
            14'h55be: o_data_a = 16'b0000000000000011;
            14'h55bf: o_data_a = 16'b1110000010100000;
            14'h55c0: o_data_a = 16'b1111110000010000;
            14'h55c1: o_data_a = 16'b0000000000000000;
            14'h55c2: o_data_a = 16'b1111110111101000;
            14'h55c3: o_data_a = 16'b1110110010100000;
            14'h55c4: o_data_a = 16'b1110001100001000;
            14'h55c5: o_data_a = 16'b0000000000000000;
            14'h55c6: o_data_a = 16'b1111110010101000;
            14'h55c7: o_data_a = 16'b1111110000010000;
            14'h55c8: o_data_a = 16'b1110110010100000;
            14'h55c9: o_data_a = 16'b1111000111001000;
            14'h55ca: o_data_a = 16'b0000000000000000;
            14'h55cb: o_data_a = 16'b1111110010101000;
            14'h55cc: o_data_a = 16'b1111110000010000;
            14'h55cd: o_data_a = 16'b0000000000000001;
            14'h55ce: o_data_a = 16'b1111110111100000;
            14'h55cf: o_data_a = 16'b1110110111100000;
            14'h55d0: o_data_a = 16'b1110110111100000;
            14'h55d1: o_data_a = 16'b1110110111100000;
            14'h55d2: o_data_a = 16'b1110110111100000;
            14'h55d3: o_data_a = 16'b1110001100001000;
            14'h55d4: o_data_a = 16'b0000000000000010;
            14'h55d5: o_data_a = 16'b1110110000010000;
            14'h55d6: o_data_a = 16'b0000000000000000;
            14'h55d7: o_data_a = 16'b1111110111101000;
            14'h55d8: o_data_a = 16'b1110110010100000;
            14'h55d9: o_data_a = 16'b1110001100001000;
            14'h55da: o_data_a = 16'b0000000000000001;
            14'h55db: o_data_a = 16'b1111110111100000;
            14'h55dc: o_data_a = 16'b1110110111100000;
            14'h55dd: o_data_a = 16'b1111110000010000;
            14'h55de: o_data_a = 16'b0000000000000000;
            14'h55df: o_data_a = 16'b1111110111101000;
            14'h55e0: o_data_a = 16'b1110110010100000;
            14'h55e1: o_data_a = 16'b1110001100001000;
            14'h55e2: o_data_a = 16'b0000000000000010;
            14'h55e3: o_data_a = 16'b1110110000010000;
            14'h55e4: o_data_a = 16'b0000000000001101;
            14'h55e5: o_data_a = 16'b1110001100001000;
            14'h55e6: o_data_a = 16'b0001101010100110;
            14'h55e7: o_data_a = 16'b1110110000010000;
            14'h55e8: o_data_a = 16'b0000000000001110;
            14'h55e9: o_data_a = 16'b1110001100001000;
            14'h55ea: o_data_a = 16'b0101010111101110;
            14'h55eb: o_data_a = 16'b1110110000010000;
            14'h55ec: o_data_a = 16'b0000000001011111;
            14'h55ed: o_data_a = 16'b1110101010000111;
            14'h55ee: o_data_a = 16'b0000000000000001;
            14'h55ef: o_data_a = 16'b1111110000010000;
            14'h55f0: o_data_a = 16'b0000000000001001;
            14'h55f1: o_data_a = 16'b1110000010010000;
            14'h55f2: o_data_a = 16'b0000000000001101;
            14'h55f3: o_data_a = 16'b1110001100001000;
            14'h55f4: o_data_a = 16'b0000000000000000;
            14'h55f5: o_data_a = 16'b1111110010101000;
            14'h55f6: o_data_a = 16'b1111110000010000;
            14'h55f7: o_data_a = 16'b0000000000001101;
            14'h55f8: o_data_a = 16'b1111110000100000;
            14'h55f9: o_data_a = 16'b1110001100001000;
            14'h55fa: o_data_a = 16'b0000000000000010;
            14'h55fb: o_data_a = 16'b1110110000010000;
            14'h55fc: o_data_a = 16'b0000000000000000;
            14'h55fd: o_data_a = 16'b1111110111101000;
            14'h55fe: o_data_a = 16'b1110110010100000;
            14'h55ff: o_data_a = 16'b1110001100001000;
            14'h5600: o_data_a = 16'b0000000000000001;
            14'h5601: o_data_a = 16'b1111110111100000;
            14'h5602: o_data_a = 16'b1110110111100000;
            14'h5603: o_data_a = 16'b1111110000010000;
            14'h5604: o_data_a = 16'b0000000000000000;
            14'h5605: o_data_a = 16'b1111110111101000;
            14'h5606: o_data_a = 16'b1110110010100000;
            14'h5607: o_data_a = 16'b1110001100001000;
            14'h5608: o_data_a = 16'b0000000000000001;
            14'h5609: o_data_a = 16'b1111110000010000;
            14'h560a: o_data_a = 16'b0000000000000011;
            14'h560b: o_data_a = 16'b1110000010100000;
            14'h560c: o_data_a = 16'b1111110000010000;
            14'h560d: o_data_a = 16'b0000000000000000;
            14'h560e: o_data_a = 16'b1111110111101000;
            14'h560f: o_data_a = 16'b1110110010100000;
            14'h5610: o_data_a = 16'b1110001100001000;
            14'h5611: o_data_a = 16'b0000000000000000;
            14'h5612: o_data_a = 16'b1111110010101000;
            14'h5613: o_data_a = 16'b1111110000010000;
            14'h5614: o_data_a = 16'b1110110010100000;
            14'h5615: o_data_a = 16'b1111000111001000;
            14'h5616: o_data_a = 16'b0000000000000010;
            14'h5617: o_data_a = 16'b1110110000010000;
            14'h5618: o_data_a = 16'b0000000000001101;
            14'h5619: o_data_a = 16'b1110001100001000;
            14'h561a: o_data_a = 16'b0001101010100110;
            14'h561b: o_data_a = 16'b1110110000010000;
            14'h561c: o_data_a = 16'b0000000000001110;
            14'h561d: o_data_a = 16'b1110001100001000;
            14'h561e: o_data_a = 16'b0101011000100010;
            14'h561f: o_data_a = 16'b1110110000010000;
            14'h5620: o_data_a = 16'b0000000001011111;
            14'h5621: o_data_a = 16'b1110101010000111;
            14'h5622: o_data_a = 16'b0000000000000001;
            14'h5623: o_data_a = 16'b1111110000010000;
            14'h5624: o_data_a = 16'b0000000000001010;
            14'h5625: o_data_a = 16'b1110000010010000;
            14'h5626: o_data_a = 16'b0000000000001101;
            14'h5627: o_data_a = 16'b1110001100001000;
            14'h5628: o_data_a = 16'b0000000000000000;
            14'h5629: o_data_a = 16'b1111110010101000;
            14'h562a: o_data_a = 16'b1111110000010000;
            14'h562b: o_data_a = 16'b0000000000001101;
            14'h562c: o_data_a = 16'b1111110000100000;
            14'h562d: o_data_a = 16'b1110001100001000;
            14'h562e: o_data_a = 16'b0000000000000001;
            14'h562f: o_data_a = 16'b1111110111100000;
            14'h5630: o_data_a = 16'b1111110000010000;
            14'h5631: o_data_a = 16'b0000000000000000;
            14'h5632: o_data_a = 16'b1111110111101000;
            14'h5633: o_data_a = 16'b1110110010100000;
            14'h5634: o_data_a = 16'b1110001100001000;
            14'h5635: o_data_a = 16'b0000000000000001;
            14'h5636: o_data_a = 16'b1111110000100000;
            14'h5637: o_data_a = 16'b1111110000010000;
            14'h5638: o_data_a = 16'b0000000000000000;
            14'h5639: o_data_a = 16'b1111110111101000;
            14'h563a: o_data_a = 16'b1110110010100000;
            14'h563b: o_data_a = 16'b1110001100001000;
            14'h563c: o_data_a = 16'b0000000000000001;
            14'h563d: o_data_a = 16'b1111110000010000;
            14'h563e: o_data_a = 16'b0000000000000110;
            14'h563f: o_data_a = 16'b1110000010100000;
            14'h5640: o_data_a = 16'b1111110000010000;
            14'h5641: o_data_a = 16'b0000000000000000;
            14'h5642: o_data_a = 16'b1111110111101000;
            14'h5643: o_data_a = 16'b1110110010100000;
            14'h5644: o_data_a = 16'b1110001100001000;
            14'h5645: o_data_a = 16'b0000000000000011;
            14'h5646: o_data_a = 16'b1110110000010000;
            14'h5647: o_data_a = 16'b0000000000001101;
            14'h5648: o_data_a = 16'b1110001100001000;
            14'h5649: o_data_a = 16'b0101001011010100;
            14'h564a: o_data_a = 16'b1110110000010000;
            14'h564b: o_data_a = 16'b0000000000001110;
            14'h564c: o_data_a = 16'b1110001100001000;
            14'h564d: o_data_a = 16'b0101011001010001;
            14'h564e: o_data_a = 16'b1110110000010000;
            14'h564f: o_data_a = 16'b0000000001011111;
            14'h5650: o_data_a = 16'b1110101010000111;
            14'h5651: o_data_a = 16'b0000000000000000;
            14'h5652: o_data_a = 16'b1111110010101000;
            14'h5653: o_data_a = 16'b1111110000010000;
            14'h5654: o_data_a = 16'b0000000000000101;
            14'h5655: o_data_a = 16'b1110001100001000;
            14'h5656: o_data_a = 16'b0000000000000001;
            14'h5657: o_data_a = 16'b1111110111100000;
            14'h5658: o_data_a = 16'b1111110000010000;
            14'h5659: o_data_a = 16'b0000000000000000;
            14'h565a: o_data_a = 16'b1111110111101000;
            14'h565b: o_data_a = 16'b1110110010100000;
            14'h565c: o_data_a = 16'b1110001100001000;
            14'h565d: o_data_a = 16'b0000000000000001;
            14'h565e: o_data_a = 16'b1111110000010000;
            14'h565f: o_data_a = 16'b0000000000001000;
            14'h5660: o_data_a = 16'b1110000010100000;
            14'h5661: o_data_a = 16'b1111110000010000;
            14'h5662: o_data_a = 16'b0000000000000000;
            14'h5663: o_data_a = 16'b1111110111101000;
            14'h5664: o_data_a = 16'b1110110010100000;
            14'h5665: o_data_a = 16'b1110001100001000;
            14'h5666: o_data_a = 16'b0101011001101010;
            14'h5667: o_data_a = 16'b1110110000010000;
            14'h5668: o_data_a = 16'b0000000000100110;
            14'h5669: o_data_a = 16'b1110101010000111;
            14'h566a: o_data_a = 16'b0000000000000000;
            14'h566b: o_data_a = 16'b1111110010100000;
            14'h566c: o_data_a = 16'b1111110001001000;
            14'h566d: o_data_a = 16'b0000000000000000;
            14'h566e: o_data_a = 16'b1111110010101000;
            14'h566f: o_data_a = 16'b1111110000010000;
            14'h5670: o_data_a = 16'b0101011101001100;
            14'h5671: o_data_a = 16'b1110001100000101;
            14'h5672: o_data_a = 16'b0000000000000001;
            14'h5673: o_data_a = 16'b1111110000010000;
            14'h5674: o_data_a = 16'b0000000000000101;
            14'h5675: o_data_a = 16'b1110000010100000;
            14'h5676: o_data_a = 16'b1111110000010000;
            14'h5677: o_data_a = 16'b0000000000000000;
            14'h5678: o_data_a = 16'b1111110111101000;
            14'h5679: o_data_a = 16'b1110110010100000;
            14'h567a: o_data_a = 16'b1110001100001000;
            14'h567b: o_data_a = 16'b0000000000000000;
            14'h567c: o_data_a = 16'b1111110111001000;
            14'h567d: o_data_a = 16'b1111110010100000;
            14'h567e: o_data_a = 16'b1110101010001000;
            14'h567f: o_data_a = 16'b0101011010000011;
            14'h5680: o_data_a = 16'b1110110000010000;
            14'h5681: o_data_a = 16'b0000000000100110;
            14'h5682: o_data_a = 16'b1110101010000111;
            14'h5683: o_data_a = 16'b0000000000000000;
            14'h5684: o_data_a = 16'b1111110010101000;
            14'h5685: o_data_a = 16'b1111110000010000;
            14'h5686: o_data_a = 16'b0101011010001010;
            14'h5687: o_data_a = 16'b1110001100000101;
            14'h5688: o_data_a = 16'b0101011010101101;
            14'h5689: o_data_a = 16'b1110101010000111;
            14'h568a: o_data_a = 16'b0000000000000001;
            14'h568b: o_data_a = 16'b1111110000010000;
            14'h568c: o_data_a = 16'b0000000000000101;
            14'h568d: o_data_a = 16'b1110000010100000;
            14'h568e: o_data_a = 16'b1111110000010000;
            14'h568f: o_data_a = 16'b0000000000000000;
            14'h5690: o_data_a = 16'b1111110111101000;
            14'h5691: o_data_a = 16'b1110110010100000;
            14'h5692: o_data_a = 16'b1110001100001000;
            14'h5693: o_data_a = 16'b0000000000000001;
            14'h5694: o_data_a = 16'b1111110000010000;
            14'h5695: o_data_a = 16'b0000000000001001;
            14'h5696: o_data_a = 16'b1110000010100000;
            14'h5697: o_data_a = 16'b1111110000010000;
            14'h5698: o_data_a = 16'b0000000000000000;
            14'h5699: o_data_a = 16'b1111110111101000;
            14'h569a: o_data_a = 16'b1110110010100000;
            14'h569b: o_data_a = 16'b1110001100001000;
            14'h569c: o_data_a = 16'b0000000000000000;
            14'h569d: o_data_a = 16'b1111110010101000;
            14'h569e: o_data_a = 16'b1111110000010000;
            14'h569f: o_data_a = 16'b1110110010100000;
            14'h56a0: o_data_a = 16'b1111000010001000;
            14'h56a1: o_data_a = 16'b0000000000000000;
            14'h56a2: o_data_a = 16'b1111110010101000;
            14'h56a3: o_data_a = 16'b1111110000010000;
            14'h56a4: o_data_a = 16'b0000000000000001;
            14'h56a5: o_data_a = 16'b1111110111100000;
            14'h56a6: o_data_a = 16'b1110110111100000;
            14'h56a7: o_data_a = 16'b1110110111100000;
            14'h56a8: o_data_a = 16'b1110110111100000;
            14'h56a9: o_data_a = 16'b1110110111100000;
            14'h56aa: o_data_a = 16'b1110001100001000;
            14'h56ab: o_data_a = 16'b0101011100001100;
            14'h56ac: o_data_a = 16'b1110101010000111;
            14'h56ad: o_data_a = 16'b0000000000000001;
            14'h56ae: o_data_a = 16'b1111110000010000;
            14'h56af: o_data_a = 16'b0000000000000101;
            14'h56b0: o_data_a = 16'b1110000010100000;
            14'h56b1: o_data_a = 16'b1111110000010000;
            14'h56b2: o_data_a = 16'b0000000000000000;
            14'h56b3: o_data_a = 16'b1111110111101000;
            14'h56b4: o_data_a = 16'b1110110010100000;
            14'h56b5: o_data_a = 16'b1110001100001000;
            14'h56b6: o_data_a = 16'b0000000000000001;
            14'h56b7: o_data_a = 16'b1111110000010000;
            14'h56b8: o_data_a = 16'b0000000000001010;
            14'h56b9: o_data_a = 16'b1110000010100000;
            14'h56ba: o_data_a = 16'b1111110000010000;
            14'h56bb: o_data_a = 16'b0000000000000000;
            14'h56bc: o_data_a = 16'b1111110111101000;
            14'h56bd: o_data_a = 16'b1110110010100000;
            14'h56be: o_data_a = 16'b1110001100001000;
            14'h56bf: o_data_a = 16'b0000000000000000;
            14'h56c0: o_data_a = 16'b1111110010101000;
            14'h56c1: o_data_a = 16'b1111110000010000;
            14'h56c2: o_data_a = 16'b1110110010100000;
            14'h56c3: o_data_a = 16'b1111000010001000;
            14'h56c4: o_data_a = 16'b0000000000000000;
            14'h56c5: o_data_a = 16'b1111110010101000;
            14'h56c6: o_data_a = 16'b1111110000010000;
            14'h56c7: o_data_a = 16'b0000000000000001;
            14'h56c8: o_data_a = 16'b1111110111100000;
            14'h56c9: o_data_a = 16'b1110110111100000;
            14'h56ca: o_data_a = 16'b1110110111100000;
            14'h56cb: o_data_a = 16'b1110110111100000;
            14'h56cc: o_data_a = 16'b1110110111100000;
            14'h56cd: o_data_a = 16'b1110001100001000;
            14'h56ce: o_data_a = 16'b0000000000000001;
            14'h56cf: o_data_a = 16'b1111110000010000;
            14'h56d0: o_data_a = 16'b0000000000000111;
            14'h56d1: o_data_a = 16'b1110000010100000;
            14'h56d2: o_data_a = 16'b1111110000010000;
            14'h56d3: o_data_a = 16'b0000000000000000;
            14'h56d4: o_data_a = 16'b1111110111101000;
            14'h56d5: o_data_a = 16'b1110110010100000;
            14'h56d6: o_data_a = 16'b1110001100001000;
            14'h56d7: o_data_a = 16'b0000000000000000;
            14'h56d8: o_data_a = 16'b1111110010101000;
            14'h56d9: o_data_a = 16'b1111110000010000;
            14'h56da: o_data_a = 16'b0101011011011110;
            14'h56db: o_data_a = 16'b1110001100000101;
            14'h56dc: o_data_a = 16'b0101011011110110;
            14'h56dd: o_data_a = 16'b1110101010000111;
            14'h56de: o_data_a = 16'b0000000000000001;
            14'h56df: o_data_a = 16'b1111110000100000;
            14'h56e0: o_data_a = 16'b1111110000010000;
            14'h56e1: o_data_a = 16'b0000000000000000;
            14'h56e2: o_data_a = 16'b1111110111101000;
            14'h56e3: o_data_a = 16'b1110110010100000;
            14'h56e4: o_data_a = 16'b1110001100001000;
            14'h56e5: o_data_a = 16'b0000000000000000;
            14'h56e6: o_data_a = 16'b1111110111001000;
            14'h56e7: o_data_a = 16'b1111110010100000;
            14'h56e8: o_data_a = 16'b1110111111001000;
            14'h56e9: o_data_a = 16'b0000000000000000;
            14'h56ea: o_data_a = 16'b1111110010101000;
            14'h56eb: o_data_a = 16'b1111110000010000;
            14'h56ec: o_data_a = 16'b1110110010100000;
            14'h56ed: o_data_a = 16'b1111000111001000;
            14'h56ee: o_data_a = 16'b0000000000000000;
            14'h56ef: o_data_a = 16'b1111110010101000;
            14'h56f0: o_data_a = 16'b1111110000010000;
            14'h56f1: o_data_a = 16'b0000000000000001;
            14'h56f2: o_data_a = 16'b1111110000100000;
            14'h56f3: o_data_a = 16'b1110001100001000;
            14'h56f4: o_data_a = 16'b0101011100001100;
            14'h56f5: o_data_a = 16'b1110101010000111;
            14'h56f6: o_data_a = 16'b0000000000000001;
            14'h56f7: o_data_a = 16'b1111110000100000;
            14'h56f8: o_data_a = 16'b1111110000010000;
            14'h56f9: o_data_a = 16'b0000000000000000;
            14'h56fa: o_data_a = 16'b1111110111101000;
            14'h56fb: o_data_a = 16'b1110110010100000;
            14'h56fc: o_data_a = 16'b1110001100001000;
            14'h56fd: o_data_a = 16'b0000000000000000;
            14'h56fe: o_data_a = 16'b1111110111001000;
            14'h56ff: o_data_a = 16'b1111110010100000;
            14'h5700: o_data_a = 16'b1110111111001000;
            14'h5701: o_data_a = 16'b0000000000000000;
            14'h5702: o_data_a = 16'b1111110010101000;
            14'h5703: o_data_a = 16'b1111110000010000;
            14'h5704: o_data_a = 16'b1110110010100000;
            14'h5705: o_data_a = 16'b1111000010001000;
            14'h5706: o_data_a = 16'b0000000000000000;
            14'h5707: o_data_a = 16'b1111110010101000;
            14'h5708: o_data_a = 16'b1111110000010000;
            14'h5709: o_data_a = 16'b0000000000000001;
            14'h570a: o_data_a = 16'b1111110000100000;
            14'h570b: o_data_a = 16'b1110001100001000;
            14'h570c: o_data_a = 16'b0000000000000001;
            14'h570d: o_data_a = 16'b1111110111100000;
            14'h570e: o_data_a = 16'b1111110000010000;
            14'h570f: o_data_a = 16'b0000000000000000;
            14'h5710: o_data_a = 16'b1111110111101000;
            14'h5711: o_data_a = 16'b1110110010100000;
            14'h5712: o_data_a = 16'b1110001100001000;
            14'h5713: o_data_a = 16'b0000000000000000;
            14'h5714: o_data_a = 16'b1111110111001000;
            14'h5715: o_data_a = 16'b1111110010100000;
            14'h5716: o_data_a = 16'b1110111111001000;
            14'h5717: o_data_a = 16'b0000000000000000;
            14'h5718: o_data_a = 16'b1111110010101000;
            14'h5719: o_data_a = 16'b1111110000010000;
            14'h571a: o_data_a = 16'b1110110010100000;
            14'h571b: o_data_a = 16'b1111000010001000;
            14'h571c: o_data_a = 16'b0000000000000000;
            14'h571d: o_data_a = 16'b1111110010101000;
            14'h571e: o_data_a = 16'b1111110000010000;
            14'h571f: o_data_a = 16'b0000000000000001;
            14'h5720: o_data_a = 16'b1111110111100000;
            14'h5721: o_data_a = 16'b1110001100001000;
            14'h5722: o_data_a = 16'b0000000000000001;
            14'h5723: o_data_a = 16'b1111110111100000;
            14'h5724: o_data_a = 16'b1111110000010000;
            14'h5725: o_data_a = 16'b0000000000000000;
            14'h5726: o_data_a = 16'b1111110111101000;
            14'h5727: o_data_a = 16'b1110110010100000;
            14'h5728: o_data_a = 16'b1110001100001000;
            14'h5729: o_data_a = 16'b0000000000000001;
            14'h572a: o_data_a = 16'b1111110000100000;
            14'h572b: o_data_a = 16'b1111110000010000;
            14'h572c: o_data_a = 16'b0000000000000000;
            14'h572d: o_data_a = 16'b1111110111101000;
            14'h572e: o_data_a = 16'b1110110010100000;
            14'h572f: o_data_a = 16'b1110001100001000;
            14'h5730: o_data_a = 16'b0000000000000001;
            14'h5731: o_data_a = 16'b1111110000010000;
            14'h5732: o_data_a = 16'b0000000000000110;
            14'h5733: o_data_a = 16'b1110000010100000;
            14'h5734: o_data_a = 16'b1111110000010000;
            14'h5735: o_data_a = 16'b0000000000000000;
            14'h5736: o_data_a = 16'b1111110111101000;
            14'h5737: o_data_a = 16'b1110110010100000;
            14'h5738: o_data_a = 16'b1110001100001000;
            14'h5739: o_data_a = 16'b0000000000000011;
            14'h573a: o_data_a = 16'b1110110000010000;
            14'h573b: o_data_a = 16'b0000000000001101;
            14'h573c: o_data_a = 16'b1110001100001000;
            14'h573d: o_data_a = 16'b0101001011010100;
            14'h573e: o_data_a = 16'b1110110000010000;
            14'h573f: o_data_a = 16'b0000000000001110;
            14'h5740: o_data_a = 16'b1110001100001000;
            14'h5741: o_data_a = 16'b0101011101000101;
            14'h5742: o_data_a = 16'b1110110000010000;
            14'h5743: o_data_a = 16'b0000000001011111;
            14'h5744: o_data_a = 16'b1110101010000111;
            14'h5745: o_data_a = 16'b0000000000000000;
            14'h5746: o_data_a = 16'b1111110010101000;
            14'h5747: o_data_a = 16'b1111110000010000;
            14'h5748: o_data_a = 16'b0000000000000101;
            14'h5749: o_data_a = 16'b1110001100001000;
            14'h574a: o_data_a = 16'b0101011001010110;
            14'h574b: o_data_a = 16'b1110101010000111;
            14'h574c: o_data_a = 16'b0000000000000000;
            14'h574d: o_data_a = 16'b1111110111001000;
            14'h574e: o_data_a = 16'b1111110010100000;
            14'h574f: o_data_a = 16'b1110101010001000;
            14'h5750: o_data_a = 16'b0000000000110110;
            14'h5751: o_data_a = 16'b1110101010000111;
            14'h5752: o_data_a = 16'b0000000000001001;
            14'h5753: o_data_a = 16'b1110110000010000;
            14'h5754: o_data_a = 16'b1110001110010000;
            14'h5755: o_data_a = 16'b0000000000000000;
            14'h5756: o_data_a = 16'b1111110111101000;
            14'h5757: o_data_a = 16'b1110110010100000;
            14'h5758: o_data_a = 16'b1110101010001000;
            14'h5759: o_data_a = 16'b0101011101010100;
            14'h575a: o_data_a = 16'b1110001100000001;
            14'h575b: o_data_a = 16'b0000000000000010;
            14'h575c: o_data_a = 16'b1111110000100000;
            14'h575d: o_data_a = 16'b1111110000010000;
            14'h575e: o_data_a = 16'b0000000000000000;
            14'h575f: o_data_a = 16'b1111110111101000;
            14'h5760: o_data_a = 16'b1110110010100000;
            14'h5761: o_data_a = 16'b1110001100001000;
            14'h5762: o_data_a = 16'b0000000000000010;
            14'h5763: o_data_a = 16'b1111110111100000;
            14'h5764: o_data_a = 16'b1110110111100000;
            14'h5765: o_data_a = 16'b1111110000010000;
            14'h5766: o_data_a = 16'b0000000000000000;
            14'h5767: o_data_a = 16'b1111110111101000;
            14'h5768: o_data_a = 16'b1110110010100000;
            14'h5769: o_data_a = 16'b1110001100001000;
            14'h576a: o_data_a = 16'b0101011101101110;
            14'h576b: o_data_a = 16'b1110110000010000;
            14'h576c: o_data_a = 16'b0000000000010110;
            14'h576d: o_data_a = 16'b1110101010000111;
            14'h576e: o_data_a = 16'b0000000000000010;
            14'h576f: o_data_a = 16'b1111110111100000;
            14'h5770: o_data_a = 16'b1111110000010000;
            14'h5771: o_data_a = 16'b0000000000000000;
            14'h5772: o_data_a = 16'b1111110111101000;
            14'h5773: o_data_a = 16'b1110110010100000;
            14'h5774: o_data_a = 16'b1110001100001000;
            14'h5775: o_data_a = 16'b0000000000000010;
            14'h5776: o_data_a = 16'b1111110000010000;
            14'h5777: o_data_a = 16'b0000000000000011;
            14'h5778: o_data_a = 16'b1110000010100000;
            14'h5779: o_data_a = 16'b1111110000010000;
            14'h577a: o_data_a = 16'b0000000000000000;
            14'h577b: o_data_a = 16'b1111110111101000;
            14'h577c: o_data_a = 16'b1110110010100000;
            14'h577d: o_data_a = 16'b1110001100001000;
            14'h577e: o_data_a = 16'b0101011110000010;
            14'h577f: o_data_a = 16'b1110110000010000;
            14'h5780: o_data_a = 16'b0000000000010110;
            14'h5781: o_data_a = 16'b1110101010000111;
            14'h5782: o_data_a = 16'b0000000000000000;
            14'h5783: o_data_a = 16'b1111110010101000;
            14'h5784: o_data_a = 16'b1111110000010000;
            14'h5785: o_data_a = 16'b1110110010100000;
            14'h5786: o_data_a = 16'b1111010101001000;
            14'h5787: o_data_a = 16'b0000000000000010;
            14'h5788: o_data_a = 16'b1111110000100000;
            14'h5789: o_data_a = 16'b1111110000010000;
            14'h578a: o_data_a = 16'b0000000000000000;
            14'h578b: o_data_a = 16'b1111110111101000;
            14'h578c: o_data_a = 16'b1110110010100000;
            14'h578d: o_data_a = 16'b1110001100001000;
            14'h578e: o_data_a = 16'b0000000000000000;
            14'h578f: o_data_a = 16'b1111110111001000;
            14'h5790: o_data_a = 16'b1111110010100000;
            14'h5791: o_data_a = 16'b1110101010001000;
            14'h5792: o_data_a = 16'b0101011110010110;
            14'h5793: o_data_a = 16'b1110110000010000;
            14'h5794: o_data_a = 16'b0000000000100110;
            14'h5795: o_data_a = 16'b1110101010000111;
            14'h5796: o_data_a = 16'b0000000000000000;
            14'h5797: o_data_a = 16'b1111110010101000;
            14'h5798: o_data_a = 16'b1111110000010000;
            14'h5799: o_data_a = 16'b1110110010100000;
            14'h579a: o_data_a = 16'b1111010101001000;
            14'h579b: o_data_a = 16'b0000000000000010;
            14'h579c: o_data_a = 16'b1111110111100000;
            14'h579d: o_data_a = 16'b1110110111100000;
            14'h579e: o_data_a = 16'b1111110000010000;
            14'h579f: o_data_a = 16'b0000000000000000;
            14'h57a0: o_data_a = 16'b1111110111101000;
            14'h57a1: o_data_a = 16'b1110110010100000;
            14'h57a2: o_data_a = 16'b1110001100001000;
            14'h57a3: o_data_a = 16'b0000000111111111;
            14'h57a4: o_data_a = 16'b1110110000010000;
            14'h57a5: o_data_a = 16'b0000000000000000;
            14'h57a6: o_data_a = 16'b1111110111101000;
            14'h57a7: o_data_a = 16'b1110110010100000;
            14'h57a8: o_data_a = 16'b1110001100001000;
            14'h57a9: o_data_a = 16'b0101011110101101;
            14'h57aa: o_data_a = 16'b1110110000010000;
            14'h57ab: o_data_a = 16'b0000000000010110;
            14'h57ac: o_data_a = 16'b1110101010000111;
            14'h57ad: o_data_a = 16'b0000000000000000;
            14'h57ae: o_data_a = 16'b1111110010101000;
            14'h57af: o_data_a = 16'b1111110000010000;
            14'h57b0: o_data_a = 16'b1110110010100000;
            14'h57b1: o_data_a = 16'b1111010101001000;
            14'h57b2: o_data_a = 16'b0000000000000010;
            14'h57b3: o_data_a = 16'b1111110111100000;
            14'h57b4: o_data_a = 16'b1111110000010000;
            14'h57b5: o_data_a = 16'b0000000000000000;
            14'h57b6: o_data_a = 16'b1111110111101000;
            14'h57b7: o_data_a = 16'b1110110010100000;
            14'h57b8: o_data_a = 16'b1110001100001000;
            14'h57b9: o_data_a = 16'b0000000000000000;
            14'h57ba: o_data_a = 16'b1111110111001000;
            14'h57bb: o_data_a = 16'b1111110010100000;
            14'h57bc: o_data_a = 16'b1110101010001000;
            14'h57bd: o_data_a = 16'b0101011111000001;
            14'h57be: o_data_a = 16'b1110110000010000;
            14'h57bf: o_data_a = 16'b0000000000100110;
            14'h57c0: o_data_a = 16'b1110101010000111;
            14'h57c1: o_data_a = 16'b0000000000000000;
            14'h57c2: o_data_a = 16'b1111110010101000;
            14'h57c3: o_data_a = 16'b1111110000010000;
            14'h57c4: o_data_a = 16'b1110110010100000;
            14'h57c5: o_data_a = 16'b1111010101001000;
            14'h57c6: o_data_a = 16'b0000000000000010;
            14'h57c7: o_data_a = 16'b1111110000010000;
            14'h57c8: o_data_a = 16'b0000000000000011;
            14'h57c9: o_data_a = 16'b1110000010100000;
            14'h57ca: o_data_a = 16'b1111110000010000;
            14'h57cb: o_data_a = 16'b0000000000000000;
            14'h57cc: o_data_a = 16'b1111110111101000;
            14'h57cd: o_data_a = 16'b1110110010100000;
            14'h57ce: o_data_a = 16'b1110001100001000;
            14'h57cf: o_data_a = 16'b0000000011111111;
            14'h57d0: o_data_a = 16'b1110110000010000;
            14'h57d1: o_data_a = 16'b0000000000000000;
            14'h57d2: o_data_a = 16'b1111110111101000;
            14'h57d3: o_data_a = 16'b1110110010100000;
            14'h57d4: o_data_a = 16'b1110001100001000;
            14'h57d5: o_data_a = 16'b0101011111011001;
            14'h57d6: o_data_a = 16'b1110110000010000;
            14'h57d7: o_data_a = 16'b0000000000010110;
            14'h57d8: o_data_a = 16'b1110101010000111;
            14'h57d9: o_data_a = 16'b0000000000000000;
            14'h57da: o_data_a = 16'b1111110010101000;
            14'h57db: o_data_a = 16'b1111110000010000;
            14'h57dc: o_data_a = 16'b1110110010100000;
            14'h57dd: o_data_a = 16'b1111010101001000;
            14'h57de: o_data_a = 16'b0000000000000000;
            14'h57df: o_data_a = 16'b1111110010101000;
            14'h57e0: o_data_a = 16'b1111110000010000;
            14'h57e1: o_data_a = 16'b0101011111100101;
            14'h57e2: o_data_a = 16'b1110001100000101;
            14'h57e3: o_data_a = 16'b0101011111111100;
            14'h57e4: o_data_a = 16'b1110101010000111;
            14'h57e5: o_data_a = 16'b0000000000001001;
            14'h57e6: o_data_a = 16'b1110110000010000;
            14'h57e7: o_data_a = 16'b0000000000000000;
            14'h57e8: o_data_a = 16'b1111110111101000;
            14'h57e9: o_data_a = 16'b1110110010100000;
            14'h57ea: o_data_a = 16'b1110001100001000;
            14'h57eb: o_data_a = 16'b0000000000000001;
            14'h57ec: o_data_a = 16'b1110110000010000;
            14'h57ed: o_data_a = 16'b0000000000001101;
            14'h57ee: o_data_a = 16'b1110001100001000;
            14'h57ef: o_data_a = 16'b0110101011011001;
            14'h57f0: o_data_a = 16'b1110110000010000;
            14'h57f1: o_data_a = 16'b0000000000001110;
            14'h57f2: o_data_a = 16'b1110001100001000;
            14'h57f3: o_data_a = 16'b0101011111110111;
            14'h57f4: o_data_a = 16'b1110110000010000;
            14'h57f5: o_data_a = 16'b0000000001011111;
            14'h57f6: o_data_a = 16'b1110101010000111;
            14'h57f7: o_data_a = 16'b0000000000000000;
            14'h57f8: o_data_a = 16'b1111110010101000;
            14'h57f9: o_data_a = 16'b1111110000010000;
            14'h57fa: o_data_a = 16'b0000000000000101;
            14'h57fb: o_data_a = 16'b1110001100001000;
            14'h57fc: o_data_a = 16'b0000000000000010;
            14'h57fd: o_data_a = 16'b1111110000100000;
            14'h57fe: o_data_a = 16'b1111110000010000;
            14'h57ff: o_data_a = 16'b0000000000000000;
            14'h5800: o_data_a = 16'b1111110111101000;
            14'h5801: o_data_a = 16'b1110110010100000;
            14'h5802: o_data_a = 16'b1110001100001000;
            14'h5803: o_data_a = 16'b0000000000010000;
            14'h5804: o_data_a = 16'b1110110000010000;
            14'h5805: o_data_a = 16'b0000000000000000;
            14'h5806: o_data_a = 16'b1111110111101000;
            14'h5807: o_data_a = 16'b1110110010100000;
            14'h5808: o_data_a = 16'b1110001100001000;
            14'h5809: o_data_a = 16'b0000000000000010;
            14'h580a: o_data_a = 16'b1110110000010000;
            14'h580b: o_data_a = 16'b0000000000001101;
            14'h580c: o_data_a = 16'b1110001100001000;
            14'h580d: o_data_a = 16'b0001110001110111;
            14'h580e: o_data_a = 16'b1110110000010000;
            14'h580f: o_data_a = 16'b0000000000001110;
            14'h5810: o_data_a = 16'b1110001100001000;
            14'h5811: o_data_a = 16'b0101100000010101;
            14'h5812: o_data_a = 16'b1110110000010000;
            14'h5813: o_data_a = 16'b0000000001011111;
            14'h5814: o_data_a = 16'b1110101010000111;
            14'h5815: o_data_a = 16'b0000000000000000;
            14'h5816: o_data_a = 16'b1111110010101000;
            14'h5817: o_data_a = 16'b1111110000010000;
            14'h5818: o_data_a = 16'b0000000000000001;
            14'h5819: o_data_a = 16'b1111110111100000;
            14'h581a: o_data_a = 16'b1110110111100000;
            14'h581b: o_data_a = 16'b1110110111100000;
            14'h581c: o_data_a = 16'b1110001100001000;
            14'h581d: o_data_a = 16'b0000000000000010;
            14'h581e: o_data_a = 16'b1111110000100000;
            14'h581f: o_data_a = 16'b1111110000010000;
            14'h5820: o_data_a = 16'b0000000000000000;
            14'h5821: o_data_a = 16'b1111110111101000;
            14'h5822: o_data_a = 16'b1110110010100000;
            14'h5823: o_data_a = 16'b1110001100001000;
            14'h5824: o_data_a = 16'b0000000000000001;
            14'h5825: o_data_a = 16'b1111110000010000;
            14'h5826: o_data_a = 16'b0000000000000011;
            14'h5827: o_data_a = 16'b1110000010100000;
            14'h5828: o_data_a = 16'b1111110000010000;
            14'h5829: o_data_a = 16'b0000000000000000;
            14'h582a: o_data_a = 16'b1111110111101000;
            14'h582b: o_data_a = 16'b1110110010100000;
            14'h582c: o_data_a = 16'b1110001100001000;
            14'h582d: o_data_a = 16'b0000000000010000;
            14'h582e: o_data_a = 16'b1110110000010000;
            14'h582f: o_data_a = 16'b0000000000000000;
            14'h5830: o_data_a = 16'b1111110111101000;
            14'h5831: o_data_a = 16'b1110110010100000;
            14'h5832: o_data_a = 16'b1110001100001000;
            14'h5833: o_data_a = 16'b0000000000000010;
            14'h5834: o_data_a = 16'b1110110000010000;
            14'h5835: o_data_a = 16'b0000000000001101;
            14'h5836: o_data_a = 16'b1110001100001000;
            14'h5837: o_data_a = 16'b0001101010100110;
            14'h5838: o_data_a = 16'b1110110000010000;
            14'h5839: o_data_a = 16'b0000000000001110;
            14'h583a: o_data_a = 16'b1110001100001000;
            14'h583b: o_data_a = 16'b0101100000111111;
            14'h583c: o_data_a = 16'b1110110000010000;
            14'h583d: o_data_a = 16'b0000000001011111;
            14'h583e: o_data_a = 16'b1110101010000111;
            14'h583f: o_data_a = 16'b0000000000000000;
            14'h5840: o_data_a = 16'b1111110010101000;
            14'h5841: o_data_a = 16'b1111110000010000;
            14'h5842: o_data_a = 16'b1110110010100000;
            14'h5843: o_data_a = 16'b1111000111001000;
            14'h5844: o_data_a = 16'b0000000000000001;
            14'h5845: o_data_a = 16'b1111110000010000;
            14'h5846: o_data_a = 16'b0000000000000111;
            14'h5847: o_data_a = 16'b1110000010010000;
            14'h5848: o_data_a = 16'b0000000000001101;
            14'h5849: o_data_a = 16'b1110001100001000;
            14'h584a: o_data_a = 16'b0000000000000000;
            14'h584b: o_data_a = 16'b1111110010101000;
            14'h584c: o_data_a = 16'b1111110000010000;
            14'h584d: o_data_a = 16'b0000000000001101;
            14'h584e: o_data_a = 16'b1111110000100000;
            14'h584f: o_data_a = 16'b1110001100001000;
            14'h5850: o_data_a = 16'b0000000000000010;
            14'h5851: o_data_a = 16'b1111110111100000;
            14'h5852: o_data_a = 16'b1110110111100000;
            14'h5853: o_data_a = 16'b1111110000010000;
            14'h5854: o_data_a = 16'b0000000000000000;
            14'h5855: o_data_a = 16'b1111110111101000;
            14'h5856: o_data_a = 16'b1110110010100000;
            14'h5857: o_data_a = 16'b1110001100001000;
            14'h5858: o_data_a = 16'b0000000000010000;
            14'h5859: o_data_a = 16'b1110110000010000;
            14'h585a: o_data_a = 16'b0000000000000000;
            14'h585b: o_data_a = 16'b1111110111101000;
            14'h585c: o_data_a = 16'b1110110010100000;
            14'h585d: o_data_a = 16'b1110001100001000;
            14'h585e: o_data_a = 16'b0000000000000010;
            14'h585f: o_data_a = 16'b1110110000010000;
            14'h5860: o_data_a = 16'b0000000000001101;
            14'h5861: o_data_a = 16'b1110001100001000;
            14'h5862: o_data_a = 16'b0001110001110111;
            14'h5863: o_data_a = 16'b1110110000010000;
            14'h5864: o_data_a = 16'b0000000000001110;
            14'h5865: o_data_a = 16'b1110001100001000;
            14'h5866: o_data_a = 16'b0101100001101010;
            14'h5867: o_data_a = 16'b1110110000010000;
            14'h5868: o_data_a = 16'b0000000001011111;
            14'h5869: o_data_a = 16'b1110101010000111;
            14'h586a: o_data_a = 16'b0000000000000000;
            14'h586b: o_data_a = 16'b1111110010101000;
            14'h586c: o_data_a = 16'b1111110000010000;
            14'h586d: o_data_a = 16'b0000000000000001;
            14'h586e: o_data_a = 16'b1111110111100000;
            14'h586f: o_data_a = 16'b1110110111100000;
            14'h5870: o_data_a = 16'b1110110111100000;
            14'h5871: o_data_a = 16'b1110110111100000;
            14'h5872: o_data_a = 16'b1110001100001000;
            14'h5873: o_data_a = 16'b0000000000000010;
            14'h5874: o_data_a = 16'b1111110111100000;
            14'h5875: o_data_a = 16'b1110110111100000;
            14'h5876: o_data_a = 16'b1111110000010000;
            14'h5877: o_data_a = 16'b0000000000000000;
            14'h5878: o_data_a = 16'b1111110111101000;
            14'h5879: o_data_a = 16'b1110110010100000;
            14'h587a: o_data_a = 16'b1110001100001000;
            14'h587b: o_data_a = 16'b0000000000000001;
            14'h587c: o_data_a = 16'b1111110000010000;
            14'h587d: o_data_a = 16'b0000000000000100;
            14'h587e: o_data_a = 16'b1110000010100000;
            14'h587f: o_data_a = 16'b1111110000010000;
            14'h5880: o_data_a = 16'b0000000000000000;
            14'h5881: o_data_a = 16'b1111110111101000;
            14'h5882: o_data_a = 16'b1110110010100000;
            14'h5883: o_data_a = 16'b1110001100001000;
            14'h5884: o_data_a = 16'b0000000000010000;
            14'h5885: o_data_a = 16'b1110110000010000;
            14'h5886: o_data_a = 16'b0000000000000000;
            14'h5887: o_data_a = 16'b1111110111101000;
            14'h5888: o_data_a = 16'b1110110010100000;
            14'h5889: o_data_a = 16'b1110001100001000;
            14'h588a: o_data_a = 16'b0000000000000010;
            14'h588b: o_data_a = 16'b1110110000010000;
            14'h588c: o_data_a = 16'b0000000000001101;
            14'h588d: o_data_a = 16'b1110001100001000;
            14'h588e: o_data_a = 16'b0001101010100110;
            14'h588f: o_data_a = 16'b1110110000010000;
            14'h5890: o_data_a = 16'b0000000000001110;
            14'h5891: o_data_a = 16'b1110001100001000;
            14'h5892: o_data_a = 16'b0101100010010110;
            14'h5893: o_data_a = 16'b1110110000010000;
            14'h5894: o_data_a = 16'b0000000001011111;
            14'h5895: o_data_a = 16'b1110101010000111;
            14'h5896: o_data_a = 16'b0000000000000000;
            14'h5897: o_data_a = 16'b1111110010101000;
            14'h5898: o_data_a = 16'b1111110000010000;
            14'h5899: o_data_a = 16'b1110110010100000;
            14'h589a: o_data_a = 16'b1111000111001000;
            14'h589b: o_data_a = 16'b0000000000000001;
            14'h589c: o_data_a = 16'b1111110000010000;
            14'h589d: o_data_a = 16'b0000000000001000;
            14'h589e: o_data_a = 16'b1110000010010000;
            14'h589f: o_data_a = 16'b0000000000001101;
            14'h58a0: o_data_a = 16'b1110001100001000;
            14'h58a1: o_data_a = 16'b0000000000000000;
            14'h58a2: o_data_a = 16'b1111110010101000;
            14'h58a3: o_data_a = 16'b1111110000010000;
            14'h58a4: o_data_a = 16'b0000000000001101;
            14'h58a5: o_data_a = 16'b1111110000100000;
            14'h58a6: o_data_a = 16'b1110001100001000;
            14'h58a7: o_data_a = 16'b0000000000000001;
            14'h58a8: o_data_a = 16'b1111110000010000;
            14'h58a9: o_data_a = 16'b0000000000000111;
            14'h58aa: o_data_a = 16'b1110000010100000;
            14'h58ab: o_data_a = 16'b1111110000010000;
            14'h58ac: o_data_a = 16'b0000000000000000;
            14'h58ad: o_data_a = 16'b1111110111101000;
            14'h58ae: o_data_a = 16'b1110110010100000;
            14'h58af: o_data_a = 16'b1110001100001000;
            14'h58b0: o_data_a = 16'b0000000000011101;
            14'h58b1: o_data_a = 16'b1111110000010000;
            14'h58b2: o_data_a = 16'b0000000000000000;
            14'h58b3: o_data_a = 16'b1111110111101000;
            14'h58b4: o_data_a = 16'b1110110010100000;
            14'h58b5: o_data_a = 16'b1110001100001000;
            14'h58b6: o_data_a = 16'b0000000000000000;
            14'h58b7: o_data_a = 16'b1111110010101000;
            14'h58b8: o_data_a = 16'b1111110000010000;
            14'h58b9: o_data_a = 16'b1110110010100000;
            14'h58ba: o_data_a = 16'b1111000010001000;
            14'h58bb: o_data_a = 16'b0000000000000000;
            14'h58bc: o_data_a = 16'b1111110010101000;
            14'h58bd: o_data_a = 16'b1111110000010000;
            14'h58be: o_data_a = 16'b0000000000000100;
            14'h58bf: o_data_a = 16'b1110001100001000;
            14'h58c0: o_data_a = 16'b0000000000000100;
            14'h58c1: o_data_a = 16'b1111110000100000;
            14'h58c2: o_data_a = 16'b1111110000010000;
            14'h58c3: o_data_a = 16'b0000000000000000;
            14'h58c4: o_data_a = 16'b1111110111101000;
            14'h58c5: o_data_a = 16'b1110110010100000;
            14'h58c6: o_data_a = 16'b1110001100001000;
            14'h58c7: o_data_a = 16'b0000000000000000;
            14'h58c8: o_data_a = 16'b1111110111001000;
            14'h58c9: o_data_a = 16'b1111110010100000;
            14'h58ca: o_data_a = 16'b1110111111001000;
            14'h58cb: o_data_a = 16'b0000000000000000;
            14'h58cc: o_data_a = 16'b1111110010101000;
            14'h58cd: o_data_a = 16'b1111110000010000;
            14'h58ce: o_data_a = 16'b1110110010100000;
            14'h58cf: o_data_a = 16'b1111000111001000;
            14'h58d0: o_data_a = 16'b0000000000000000;
            14'h58d1: o_data_a = 16'b1111110010100000;
            14'h58d2: o_data_a = 16'b1111110001001000;
            14'h58d3: o_data_a = 16'b0000000000000000;
            14'h58d4: o_data_a = 16'b1111110010101000;
            14'h58d5: o_data_a = 16'b1111110000010000;
            14'h58d6: o_data_a = 16'b0000000000000001;
            14'h58d7: o_data_a = 16'b1111110111100000;
            14'h58d8: o_data_a = 16'b1110110111100000;
            14'h58d9: o_data_a = 16'b1110110111100000;
            14'h58da: o_data_a = 16'b1110110111100000;
            14'h58db: o_data_a = 16'b1110110111100000;
            14'h58dc: o_data_a = 16'b1110110111100000;
            14'h58dd: o_data_a = 16'b1110001100001000;
            14'h58de: o_data_a = 16'b0000000000000001;
            14'h58df: o_data_a = 16'b1111110000010000;
            14'h58e0: o_data_a = 16'b0000000000001000;
            14'h58e1: o_data_a = 16'b1110000010100000;
            14'h58e2: o_data_a = 16'b1111110000010000;
            14'h58e3: o_data_a = 16'b0000000000000000;
            14'h58e4: o_data_a = 16'b1111110111101000;
            14'h58e5: o_data_a = 16'b1110110010100000;
            14'h58e6: o_data_a = 16'b1110001100001000;
            14'h58e7: o_data_a = 16'b0000000000000000;
            14'h58e8: o_data_a = 16'b1111110111001000;
            14'h58e9: o_data_a = 16'b1111110010100000;
            14'h58ea: o_data_a = 16'b1110111111001000;
            14'h58eb: o_data_a = 16'b0000000000000000;
            14'h58ec: o_data_a = 16'b1111110010101000;
            14'h58ed: o_data_a = 16'b1111110000010000;
            14'h58ee: o_data_a = 16'b1110110010100000;
            14'h58ef: o_data_a = 16'b1111000010001000;
            14'h58f0: o_data_a = 16'b0000000000011101;
            14'h58f1: o_data_a = 16'b1111110000010000;
            14'h58f2: o_data_a = 16'b0000000000000000;
            14'h58f3: o_data_a = 16'b1111110111101000;
            14'h58f4: o_data_a = 16'b1110110010100000;
            14'h58f5: o_data_a = 16'b1110001100001000;
            14'h58f6: o_data_a = 16'b0000000000000000;
            14'h58f7: o_data_a = 16'b1111110010101000;
            14'h58f8: o_data_a = 16'b1111110000010000;
            14'h58f9: o_data_a = 16'b1110110010100000;
            14'h58fa: o_data_a = 16'b1111000010001000;
            14'h58fb: o_data_a = 16'b0000000000000000;
            14'h58fc: o_data_a = 16'b1111110010101000;
            14'h58fd: o_data_a = 16'b1111110000010000;
            14'h58fe: o_data_a = 16'b0000000000000100;
            14'h58ff: o_data_a = 16'b1110001100001000;
            14'h5900: o_data_a = 16'b0000000000000100;
            14'h5901: o_data_a = 16'b1111110000100000;
            14'h5902: o_data_a = 16'b1111110000010000;
            14'h5903: o_data_a = 16'b0000000000000000;
            14'h5904: o_data_a = 16'b1111110111101000;
            14'h5905: o_data_a = 16'b1110110010100000;
            14'h5906: o_data_a = 16'b1110001100001000;
            14'h5907: o_data_a = 16'b0000000000000000;
            14'h5908: o_data_a = 16'b1111110111001000;
            14'h5909: o_data_a = 16'b1111110010100000;
            14'h590a: o_data_a = 16'b1110111111001000;
            14'h590b: o_data_a = 16'b0000000000000000;
            14'h590c: o_data_a = 16'b1111110010101000;
            14'h590d: o_data_a = 16'b1111110000010000;
            14'h590e: o_data_a = 16'b1110110010100000;
            14'h590f: o_data_a = 16'b1111000111001000;
            14'h5910: o_data_a = 16'b0000000000000000;
            14'h5911: o_data_a = 16'b1111110010101000;
            14'h5912: o_data_a = 16'b1111110000010000;
            14'h5913: o_data_a = 16'b0000000000000001;
            14'h5914: o_data_a = 16'b1111110111100000;
            14'h5915: o_data_a = 16'b1110110111100000;
            14'h5916: o_data_a = 16'b1110110111100000;
            14'h5917: o_data_a = 16'b1110110111100000;
            14'h5918: o_data_a = 16'b1110110111100000;
            14'h5919: o_data_a = 16'b1110001100001000;
            14'h591a: o_data_a = 16'b0000000000000010;
            14'h591b: o_data_a = 16'b1111110111100000;
            14'h591c: o_data_a = 16'b1111110000010000;
            14'h591d: o_data_a = 16'b0000000000000000;
            14'h591e: o_data_a = 16'b1111110111101000;
            14'h591f: o_data_a = 16'b1110110010100000;
            14'h5920: o_data_a = 16'b1110001100001000;
            14'h5921: o_data_a = 16'b0000000000100000;
            14'h5922: o_data_a = 16'b1110110000010000;
            14'h5923: o_data_a = 16'b0000000000000000;
            14'h5924: o_data_a = 16'b1111110111101000;
            14'h5925: o_data_a = 16'b1110110010100000;
            14'h5926: o_data_a = 16'b1110001100001000;
            14'h5927: o_data_a = 16'b0000000000000010;
            14'h5928: o_data_a = 16'b1110110000010000;
            14'h5929: o_data_a = 16'b0000000000001101;
            14'h592a: o_data_a = 16'b1110001100001000;
            14'h592b: o_data_a = 16'b0001101010100110;
            14'h592c: o_data_a = 16'b1110110000010000;
            14'h592d: o_data_a = 16'b0000000000001110;
            14'h592e: o_data_a = 16'b1110001100001000;
            14'h592f: o_data_a = 16'b0101100100110011;
            14'h5930: o_data_a = 16'b1110110000010000;
            14'h5931: o_data_a = 16'b0000000001011111;
            14'h5932: o_data_a = 16'b1110101010000111;
            14'h5933: o_data_a = 16'b0000000000000001;
            14'h5934: o_data_a = 16'b1111110000010000;
            14'h5935: o_data_a = 16'b0000000000000011;
            14'h5936: o_data_a = 16'b1110000010100000;
            14'h5937: o_data_a = 16'b1111110000010000;
            14'h5938: o_data_a = 16'b0000000000000000;
            14'h5939: o_data_a = 16'b1111110111101000;
            14'h593a: o_data_a = 16'b1110110010100000;
            14'h593b: o_data_a = 16'b1110001100001000;
            14'h593c: o_data_a = 16'b0000000000000000;
            14'h593d: o_data_a = 16'b1111110010101000;
            14'h593e: o_data_a = 16'b1111110000010000;
            14'h593f: o_data_a = 16'b1110110010100000;
            14'h5940: o_data_a = 16'b1111000010001000;
            14'h5941: o_data_a = 16'b0000000000000000;
            14'h5942: o_data_a = 16'b1111110010101000;
            14'h5943: o_data_a = 16'b1111110000010000;
            14'h5944: o_data_a = 16'b0000000000000001;
            14'h5945: o_data_a = 16'b1111110000100000;
            14'h5946: o_data_a = 16'b1110001100001000;
            14'h5947: o_data_a = 16'b0000000000000001;
            14'h5948: o_data_a = 16'b1111110000010000;
            14'h5949: o_data_a = 16'b0000000000000100;
            14'h594a: o_data_a = 16'b1110000010100000;
            14'h594b: o_data_a = 16'b1111110000010000;
            14'h594c: o_data_a = 16'b0000000000000000;
            14'h594d: o_data_a = 16'b1111110111101000;
            14'h594e: o_data_a = 16'b1110110010100000;
            14'h594f: o_data_a = 16'b1110001100001000;
            14'h5950: o_data_a = 16'b0000000000000001;
            14'h5951: o_data_a = 16'b1111110000010000;
            14'h5952: o_data_a = 16'b0000000000000011;
            14'h5953: o_data_a = 16'b1110000010100000;
            14'h5954: o_data_a = 16'b1111110000010000;
            14'h5955: o_data_a = 16'b0000000000000000;
            14'h5956: o_data_a = 16'b1111110111101000;
            14'h5957: o_data_a = 16'b1110110010100000;
            14'h5958: o_data_a = 16'b1110001100001000;
            14'h5959: o_data_a = 16'b0000000000000000;
            14'h595a: o_data_a = 16'b1111110010101000;
            14'h595b: o_data_a = 16'b1111110000010000;
            14'h595c: o_data_a = 16'b1110110010100000;
            14'h595d: o_data_a = 16'b1111000111001000;
            14'h595e: o_data_a = 16'b0000000000000000;
            14'h595f: o_data_a = 16'b1111110010101000;
            14'h5960: o_data_a = 16'b1111110000010000;
            14'h5961: o_data_a = 16'b0000000000000001;
            14'h5962: o_data_a = 16'b1111110111100000;
            14'h5963: o_data_a = 16'b1110110111100000;
            14'h5964: o_data_a = 16'b1110001100001000;
            14'h5965: o_data_a = 16'b0000000000000010;
            14'h5966: o_data_a = 16'b1111110111100000;
            14'h5967: o_data_a = 16'b1111110000010000;
            14'h5968: o_data_a = 16'b0000000000000000;
            14'h5969: o_data_a = 16'b1111110111101000;
            14'h596a: o_data_a = 16'b1110110010100000;
            14'h596b: o_data_a = 16'b1110001100001000;
            14'h596c: o_data_a = 16'b0000000000000010;
            14'h596d: o_data_a = 16'b1111110000010000;
            14'h596e: o_data_a = 16'b0000000000000011;
            14'h596f: o_data_a = 16'b1110000010100000;
            14'h5970: o_data_a = 16'b1111110000010000;
            14'h5971: o_data_a = 16'b0000000000000000;
            14'h5972: o_data_a = 16'b1111110111101000;
            14'h5973: o_data_a = 16'b1110110010100000;
            14'h5974: o_data_a = 16'b1110001100001000;
            14'h5975: o_data_a = 16'b0101100101111001;
            14'h5976: o_data_a = 16'b1110110000010000;
            14'h5977: o_data_a = 16'b0000000000010110;
            14'h5978: o_data_a = 16'b1110101010000111;
            14'h5979: o_data_a = 16'b0000000000000000;
            14'h597a: o_data_a = 16'b1111110010100000;
            14'h597b: o_data_a = 16'b1111110001001000;
            14'h597c: o_data_a = 16'b0000000000000000;
            14'h597d: o_data_a = 16'b1111110010100000;
            14'h597e: o_data_a = 16'b1111110001001000;
            14'h597f: o_data_a = 16'b0000000000000000;
            14'h5980: o_data_a = 16'b1111110010101000;
            14'h5981: o_data_a = 16'b1111110000010000;
            14'h5982: o_data_a = 16'b0101101011001101;
            14'h5983: o_data_a = 16'b1110001100000101;
            14'h5984: o_data_a = 16'b0000000000000001;
            14'h5985: o_data_a = 16'b1111110000100000;
            14'h5986: o_data_a = 16'b1111110000010000;
            14'h5987: o_data_a = 16'b0000000000000000;
            14'h5988: o_data_a = 16'b1111110111101000;
            14'h5989: o_data_a = 16'b1110110010100000;
            14'h598a: o_data_a = 16'b1110001100001000;
            14'h598b: o_data_a = 16'b0000000000000001;
            14'h598c: o_data_a = 16'b1111110111100000;
            14'h598d: o_data_a = 16'b1110110111100000;
            14'h598e: o_data_a = 16'b1111110000010000;
            14'h598f: o_data_a = 16'b0000000000000000;
            14'h5990: o_data_a = 16'b1111110111101000;
            14'h5991: o_data_a = 16'b1110110010100000;
            14'h5992: o_data_a = 16'b1110001100001000;
            14'h5993: o_data_a = 16'b0000000000000000;
            14'h5994: o_data_a = 16'b1111110010101000;
            14'h5995: o_data_a = 16'b1111110000010000;
            14'h5996: o_data_a = 16'b1110110010100000;
            14'h5997: o_data_a = 16'b1111000010001000;
            14'h5998: o_data_a = 16'b0000000000000000;
            14'h5999: o_data_a = 16'b1111110010101000;
            14'h599a: o_data_a = 16'b1111110000010000;
            14'h599b: o_data_a = 16'b0000000000000001;
            14'h599c: o_data_a = 16'b1111110111100000;
            14'h599d: o_data_a = 16'b1110001100001000;
            14'h599e: o_data_a = 16'b0000000000000001;
            14'h599f: o_data_a = 16'b1111110111100000;
            14'h59a0: o_data_a = 16'b1110110111100000;
            14'h59a1: o_data_a = 16'b1111110000010000;
            14'h59a2: o_data_a = 16'b0000000000000000;
            14'h59a3: o_data_a = 16'b1111110111101000;
            14'h59a4: o_data_a = 16'b1110110010100000;
            14'h59a5: o_data_a = 16'b1110001100001000;
            14'h59a6: o_data_a = 16'b0000000000000000;
            14'h59a7: o_data_a = 16'b1111110111001000;
            14'h59a8: o_data_a = 16'b1111110010100000;
            14'h59a9: o_data_a = 16'b1110101010001000;
            14'h59aa: o_data_a = 16'b0101100110101110;
            14'h59ab: o_data_a = 16'b1110110000010000;
            14'h59ac: o_data_a = 16'b0000000000000110;
            14'h59ad: o_data_a = 16'b1110101010000111;
            14'h59ae: o_data_a = 16'b0000000000000000;
            14'h59af: o_data_a = 16'b1111110010101000;
            14'h59b0: o_data_a = 16'b1111110000010000;
            14'h59b1: o_data_a = 16'b0101100110110101;
            14'h59b2: o_data_a = 16'b1110001100000101;
            14'h59b3: o_data_a = 16'b0101100111100110;
            14'h59b4: o_data_a = 16'b1110101010000111;
            14'h59b5: o_data_a = 16'b0000000000000001;
            14'h59b6: o_data_a = 16'b1111110000100000;
            14'h59b7: o_data_a = 16'b1111110000010000;
            14'h59b8: o_data_a = 16'b0000000000000000;
            14'h59b9: o_data_a = 16'b1111110111101000;
            14'h59ba: o_data_a = 16'b1110110010100000;
            14'h59bb: o_data_a = 16'b1110001100001000;
            14'h59bc: o_data_a = 16'b0000000000000001;
            14'h59bd: o_data_a = 16'b1111110000010000;
            14'h59be: o_data_a = 16'b0000000000000101;
            14'h59bf: o_data_a = 16'b1110000010100000;
            14'h59c0: o_data_a = 16'b1111110000010000;
            14'h59c1: o_data_a = 16'b0000000000000000;
            14'h59c2: o_data_a = 16'b1111110111101000;
            14'h59c3: o_data_a = 16'b1110110010100000;
            14'h59c4: o_data_a = 16'b1110001100001000;
            14'h59c5: o_data_a = 16'b0000000000000001;
            14'h59c6: o_data_a = 16'b1111110000010000;
            14'h59c7: o_data_a = 16'b0000000000000110;
            14'h59c8: o_data_a = 16'b1110000010100000;
            14'h59c9: o_data_a = 16'b1111110000010000;
            14'h59ca: o_data_a = 16'b0000000000000000;
            14'h59cb: o_data_a = 16'b1111110111101000;
            14'h59cc: o_data_a = 16'b1110110010100000;
            14'h59cd: o_data_a = 16'b1110001100001000;
            14'h59ce: o_data_a = 16'b0000000000000000;
            14'h59cf: o_data_a = 16'b1111110010101000;
            14'h59d0: o_data_a = 16'b1111110000010000;
            14'h59d1: o_data_a = 16'b1110110010100000;
            14'h59d2: o_data_a = 16'b1111000000001000;
            14'h59d3: o_data_a = 16'b0000000000000010;
            14'h59d4: o_data_a = 16'b1110110000010000;
            14'h59d5: o_data_a = 16'b0000000000001101;
            14'h59d6: o_data_a = 16'b1110001100001000;
            14'h59d7: o_data_a = 16'b0101000011011101;
            14'h59d8: o_data_a = 16'b1110110000010000;
            14'h59d9: o_data_a = 16'b0000000000001110;
            14'h59da: o_data_a = 16'b1110001100001000;
            14'h59db: o_data_a = 16'b0101100111011111;
            14'h59dc: o_data_a = 16'b1110110000010000;
            14'h59dd: o_data_a = 16'b0000000001011111;
            14'h59de: o_data_a = 16'b1110101010000111;
            14'h59df: o_data_a = 16'b0000000000000000;
            14'h59e0: o_data_a = 16'b1111110010101000;
            14'h59e1: o_data_a = 16'b1111110000010000;
            14'h59e2: o_data_a = 16'b0000000000000101;
            14'h59e3: o_data_a = 16'b1110001100001000;
            14'h59e4: o_data_a = 16'b0101101010010000;
            14'h59e5: o_data_a = 16'b1110101010000111;
            14'h59e6: o_data_a = 16'b0000000000000001;
            14'h59e7: o_data_a = 16'b1111110000100000;
            14'h59e8: o_data_a = 16'b1111110000010000;
            14'h59e9: o_data_a = 16'b0000000000000000;
            14'h59ea: o_data_a = 16'b1111110111101000;
            14'h59eb: o_data_a = 16'b1110110010100000;
            14'h59ec: o_data_a = 16'b1110001100001000;
            14'h59ed: o_data_a = 16'b0000000000000001;
            14'h59ee: o_data_a = 16'b1111110000010000;
            14'h59ef: o_data_a = 16'b0000000000000110;
            14'h59f0: o_data_a = 16'b1110000010100000;
            14'h59f1: o_data_a = 16'b1111110000010000;
            14'h59f2: o_data_a = 16'b0000000000000000;
            14'h59f3: o_data_a = 16'b1111110111101000;
            14'h59f4: o_data_a = 16'b1110110010100000;
            14'h59f5: o_data_a = 16'b1110001100001000;
            14'h59f6: o_data_a = 16'b0000000000000010;
            14'h59f7: o_data_a = 16'b1110110000010000;
            14'h59f8: o_data_a = 16'b0000000000001101;
            14'h59f9: o_data_a = 16'b1110001100001000;
            14'h59fa: o_data_a = 16'b0101000011011101;
            14'h59fb: o_data_a = 16'b1110110000010000;
            14'h59fc: o_data_a = 16'b0000000000001110;
            14'h59fd: o_data_a = 16'b1110001100001000;
            14'h59fe: o_data_a = 16'b0101101000000010;
            14'h59ff: o_data_a = 16'b1110110000010000;
            14'h5a00: o_data_a = 16'b0000000001011111;
            14'h5a01: o_data_a = 16'b1110101010000111;
            14'h5a02: o_data_a = 16'b0000000000000000;
            14'h5a03: o_data_a = 16'b1111110010101000;
            14'h5a04: o_data_a = 16'b1111110000010000;
            14'h5a05: o_data_a = 16'b0000000000000101;
            14'h5a06: o_data_a = 16'b1110001100001000;
            14'h5a07: o_data_a = 16'b0000000000000001;
            14'h5a08: o_data_a = 16'b1111110000100000;
            14'h5a09: o_data_a = 16'b1111110000010000;
            14'h5a0a: o_data_a = 16'b0000000000000000;
            14'h5a0b: o_data_a = 16'b1111110111101000;
            14'h5a0c: o_data_a = 16'b1110110010100000;
            14'h5a0d: o_data_a = 16'b1110001100001000;
            14'h5a0e: o_data_a = 16'b0000000000000000;
            14'h5a0f: o_data_a = 16'b1111110111001000;
            14'h5a10: o_data_a = 16'b1111110010100000;
            14'h5a11: o_data_a = 16'b1110111111001000;
            14'h5a12: o_data_a = 16'b0000000000000000;
            14'h5a13: o_data_a = 16'b1111110010101000;
            14'h5a14: o_data_a = 16'b1111110000010000;
            14'h5a15: o_data_a = 16'b1110110010100000;
            14'h5a16: o_data_a = 16'b1111000010001000;
            14'h5a17: o_data_a = 16'b0000000000000000;
            14'h5a18: o_data_a = 16'b1111110010101000;
            14'h5a19: o_data_a = 16'b1111110000010000;
            14'h5a1a: o_data_a = 16'b0000000000000001;
            14'h5a1b: o_data_a = 16'b1111110000100000;
            14'h5a1c: o_data_a = 16'b1110001100001000;
            14'h5a1d: o_data_a = 16'b0000000000000001;
            14'h5a1e: o_data_a = 16'b1111110000100000;
            14'h5a1f: o_data_a = 16'b1111110000010000;
            14'h5a20: o_data_a = 16'b0000000000000000;
            14'h5a21: o_data_a = 16'b1111110111101000;
            14'h5a22: o_data_a = 16'b1110110010100000;
            14'h5a23: o_data_a = 16'b1110001100001000;
            14'h5a24: o_data_a = 16'b0000000000000001;
            14'h5a25: o_data_a = 16'b1111110111100000;
            14'h5a26: o_data_a = 16'b1111110000010000;
            14'h5a27: o_data_a = 16'b0000000000000000;
            14'h5a28: o_data_a = 16'b1111110111101000;
            14'h5a29: o_data_a = 16'b1110110010100000;
            14'h5a2a: o_data_a = 16'b1110001100001000;
            14'h5a2b: o_data_a = 16'b0101101000101111;
            14'h5a2c: o_data_a = 16'b1110110000010000;
            14'h5a2d: o_data_a = 16'b0000000000100110;
            14'h5a2e: o_data_a = 16'b1110101010000111;
            14'h5a2f: o_data_a = 16'b0000000000000000;
            14'h5a30: o_data_a = 16'b1111110010100000;
            14'h5a31: o_data_a = 16'b1111110001001000;
            14'h5a32: o_data_a = 16'b0000000000000000;
            14'h5a33: o_data_a = 16'b1111110010101000;
            14'h5a34: o_data_a = 16'b1111110000010000;
            14'h5a35: o_data_a = 16'b0101101001101111;
            14'h5a36: o_data_a = 16'b1110001100000101;
            14'h5a37: o_data_a = 16'b0000000000000001;
            14'h5a38: o_data_a = 16'b1111110000100000;
            14'h5a39: o_data_a = 16'b1111110000010000;
            14'h5a3a: o_data_a = 16'b0000000000000000;
            14'h5a3b: o_data_a = 16'b1111110111101000;
            14'h5a3c: o_data_a = 16'b1110110010100000;
            14'h5a3d: o_data_a = 16'b1110001100001000;
            14'h5a3e: o_data_a = 16'b0000000000000000;
            14'h5a3f: o_data_a = 16'b1111110111001000;
            14'h5a40: o_data_a = 16'b1111110010100000;
            14'h5a41: o_data_a = 16'b1110111111001000;
            14'h5a42: o_data_a = 16'b0000000000000000;
            14'h5a43: o_data_a = 16'b1111110010100000;
            14'h5a44: o_data_a = 16'b1111110001010000;
            14'h5a45: o_data_a = 16'b1110011111001000;
            14'h5a46: o_data_a = 16'b0000000000000010;
            14'h5a47: o_data_a = 16'b1110110000010000;
            14'h5a48: o_data_a = 16'b0000000000001101;
            14'h5a49: o_data_a = 16'b1110001100001000;
            14'h5a4a: o_data_a = 16'b0101000011011101;
            14'h5a4b: o_data_a = 16'b1110110000010000;
            14'h5a4c: o_data_a = 16'b0000000000001110;
            14'h5a4d: o_data_a = 16'b1110001100001000;
            14'h5a4e: o_data_a = 16'b0101101001010010;
            14'h5a4f: o_data_a = 16'b1110110000010000;
            14'h5a50: o_data_a = 16'b0000000001011111;
            14'h5a51: o_data_a = 16'b1110101010000111;
            14'h5a52: o_data_a = 16'b0000000000000000;
            14'h5a53: o_data_a = 16'b1111110010101000;
            14'h5a54: o_data_a = 16'b1111110000010000;
            14'h5a55: o_data_a = 16'b0000000000000101;
            14'h5a56: o_data_a = 16'b1110001100001000;
            14'h5a57: o_data_a = 16'b0000000000000001;
            14'h5a58: o_data_a = 16'b1111110000100000;
            14'h5a59: o_data_a = 16'b1111110000010000;
            14'h5a5a: o_data_a = 16'b0000000000000000;
            14'h5a5b: o_data_a = 16'b1111110111101000;
            14'h5a5c: o_data_a = 16'b1110110010100000;
            14'h5a5d: o_data_a = 16'b1110001100001000;
            14'h5a5e: o_data_a = 16'b0000000000000000;
            14'h5a5f: o_data_a = 16'b1111110111001000;
            14'h5a60: o_data_a = 16'b1111110010100000;
            14'h5a61: o_data_a = 16'b1110111111001000;
            14'h5a62: o_data_a = 16'b0000000000000000;
            14'h5a63: o_data_a = 16'b1111110010101000;
            14'h5a64: o_data_a = 16'b1111110000010000;
            14'h5a65: o_data_a = 16'b1110110010100000;
            14'h5a66: o_data_a = 16'b1111000010001000;
            14'h5a67: o_data_a = 16'b0000000000000000;
            14'h5a68: o_data_a = 16'b1111110010101000;
            14'h5a69: o_data_a = 16'b1111110000010000;
            14'h5a6a: o_data_a = 16'b0000000000000001;
            14'h5a6b: o_data_a = 16'b1111110000100000;
            14'h5a6c: o_data_a = 16'b1110001100001000;
            14'h5a6d: o_data_a = 16'b0101101000011101;
            14'h5a6e: o_data_a = 16'b1110101010000111;
            14'h5a6f: o_data_a = 16'b0000000000000001;
            14'h5a70: o_data_a = 16'b1111110111100000;
            14'h5a71: o_data_a = 16'b1111110000010000;
            14'h5a72: o_data_a = 16'b0000000000000000;
            14'h5a73: o_data_a = 16'b1111110111101000;
            14'h5a74: o_data_a = 16'b1110110010100000;
            14'h5a75: o_data_a = 16'b1110001100001000;
            14'h5a76: o_data_a = 16'b0000000000000001;
            14'h5a77: o_data_a = 16'b1111110000010000;
            14'h5a78: o_data_a = 16'b0000000000000101;
            14'h5a79: o_data_a = 16'b1110000010100000;
            14'h5a7a: o_data_a = 16'b1111110000010000;
            14'h5a7b: o_data_a = 16'b0000000000000000;
            14'h5a7c: o_data_a = 16'b1111110111101000;
            14'h5a7d: o_data_a = 16'b1110110010100000;
            14'h5a7e: o_data_a = 16'b1110001100001000;
            14'h5a7f: o_data_a = 16'b0000000000000010;
            14'h5a80: o_data_a = 16'b1110110000010000;
            14'h5a81: o_data_a = 16'b0000000000001101;
            14'h5a82: o_data_a = 16'b1110001100001000;
            14'h5a83: o_data_a = 16'b0101000011011101;
            14'h5a84: o_data_a = 16'b1110110000010000;
            14'h5a85: o_data_a = 16'b0000000000001110;
            14'h5a86: o_data_a = 16'b1110001100001000;
            14'h5a87: o_data_a = 16'b0101101010001011;
            14'h5a88: o_data_a = 16'b1110110000010000;
            14'h5a89: o_data_a = 16'b0000000001011111;
            14'h5a8a: o_data_a = 16'b1110101010000111;
            14'h5a8b: o_data_a = 16'b0000000000000000;
            14'h5a8c: o_data_a = 16'b1111110010101000;
            14'h5a8d: o_data_a = 16'b1111110000010000;
            14'h5a8e: o_data_a = 16'b0000000000000101;
            14'h5a8f: o_data_a = 16'b1110001100001000;
            14'h5a90: o_data_a = 16'b0000000000000010;
            14'h5a91: o_data_a = 16'b1111110111100000;
            14'h5a92: o_data_a = 16'b1111110000010000;
            14'h5a93: o_data_a = 16'b0000000000000000;
            14'h5a94: o_data_a = 16'b1111110111101000;
            14'h5a95: o_data_a = 16'b1110110010100000;
            14'h5a96: o_data_a = 16'b1110001100001000;
            14'h5a97: o_data_a = 16'b0000000000000000;
            14'h5a98: o_data_a = 16'b1111110111001000;
            14'h5a99: o_data_a = 16'b1111110010100000;
            14'h5a9a: o_data_a = 16'b1110111111001000;
            14'h5a9b: o_data_a = 16'b0000000000000000;
            14'h5a9c: o_data_a = 16'b1111110010101000;
            14'h5a9d: o_data_a = 16'b1111110000010000;
            14'h5a9e: o_data_a = 16'b1110110010100000;
            14'h5a9f: o_data_a = 16'b1111000010001000;
            14'h5aa0: o_data_a = 16'b0000000000000000;
            14'h5aa1: o_data_a = 16'b1111110010101000;
            14'h5aa2: o_data_a = 16'b1111110000010000;
            14'h5aa3: o_data_a = 16'b0000000000000010;
            14'h5aa4: o_data_a = 16'b1111110111100000;
            14'h5aa5: o_data_a = 16'b1110001100001000;
            14'h5aa6: o_data_a = 16'b0000000000000001;
            14'h5aa7: o_data_a = 16'b1111110111100000;
            14'h5aa8: o_data_a = 16'b1111110000010000;
            14'h5aa9: o_data_a = 16'b0000000000000000;
            14'h5aaa: o_data_a = 16'b1111110111101000;
            14'h5aab: o_data_a = 16'b1110110010100000;
            14'h5aac: o_data_a = 16'b1110001100001000;
            14'h5aad: o_data_a = 16'b0000000000100000;
            14'h5aae: o_data_a = 16'b1110110000010000;
            14'h5aaf: o_data_a = 16'b0000000000000000;
            14'h5ab0: o_data_a = 16'b1111110111101000;
            14'h5ab1: o_data_a = 16'b1110110010100000;
            14'h5ab2: o_data_a = 16'b1110001100001000;
            14'h5ab3: o_data_a = 16'b0000000000000000;
            14'h5ab4: o_data_a = 16'b1111110010101000;
            14'h5ab5: o_data_a = 16'b1111110000010000;
            14'h5ab6: o_data_a = 16'b1110110010100000;
            14'h5ab7: o_data_a = 16'b1111000010001000;
            14'h5ab8: o_data_a = 16'b0000000000000001;
            14'h5ab9: o_data_a = 16'b1111110111100000;
            14'h5aba: o_data_a = 16'b1110110111100000;
            14'h5abb: o_data_a = 16'b1111110000010000;
            14'h5abc: o_data_a = 16'b0000000000000000;
            14'h5abd: o_data_a = 16'b1111110111101000;
            14'h5abe: o_data_a = 16'b1110110010100000;
            14'h5abf: o_data_a = 16'b1110001100001000;
            14'h5ac0: o_data_a = 16'b0000000000000000;
            14'h5ac1: o_data_a = 16'b1111110010101000;
            14'h5ac2: o_data_a = 16'b1111110000010000;
            14'h5ac3: o_data_a = 16'b1110110010100000;
            14'h5ac4: o_data_a = 16'b1111000111001000;
            14'h5ac5: o_data_a = 16'b0000000000000000;
            14'h5ac6: o_data_a = 16'b1111110010101000;
            14'h5ac7: o_data_a = 16'b1111110000010000;
            14'h5ac8: o_data_a = 16'b0000000000000001;
            14'h5ac9: o_data_a = 16'b1111110000100000;
            14'h5aca: o_data_a = 16'b1110001100001000;
            14'h5acb: o_data_a = 16'b0101100101100101;
            14'h5acc: o_data_a = 16'b1110101010000111;
            14'h5acd: o_data_a = 16'b0000000000000000;
            14'h5ace: o_data_a = 16'b1111110111001000;
            14'h5acf: o_data_a = 16'b1111110010100000;
            14'h5ad0: o_data_a = 16'b1110101010001000;
            14'h5ad1: o_data_a = 16'b0000000000110110;
            14'h5ad2: o_data_a = 16'b1110101010000111;
            14'h5ad3: o_data_a = 16'b0000000000001011;
            14'h5ad4: o_data_a = 16'b1110110000010000;
            14'h5ad5: o_data_a = 16'b1110001110010000;
            14'h5ad6: o_data_a = 16'b0000000000000000;
            14'h5ad7: o_data_a = 16'b1111110111101000;
            14'h5ad8: o_data_a = 16'b1110110010100000;
            14'h5ad9: o_data_a = 16'b1110101010001000;
            14'h5ada: o_data_a = 16'b0101101011010101;
            14'h5adb: o_data_a = 16'b1110001100000001;
            14'h5adc: o_data_a = 16'b0000000000000010;
            14'h5add: o_data_a = 16'b1111110111100000;
            14'h5ade: o_data_a = 16'b1111110000010000;
            14'h5adf: o_data_a = 16'b0000000000000000;
            14'h5ae0: o_data_a = 16'b1111110111101000;
            14'h5ae1: o_data_a = 16'b1110110010100000;
            14'h5ae2: o_data_a = 16'b1110001100001000;
            14'h5ae3: o_data_a = 16'b0000000000000010;
            14'h5ae4: o_data_a = 16'b1111110111100000;
            14'h5ae5: o_data_a = 16'b1110110111100000;
            14'h5ae6: o_data_a = 16'b1111110000010000;
            14'h5ae7: o_data_a = 16'b0000000000000000;
            14'h5ae8: o_data_a = 16'b1111110111101000;
            14'h5ae9: o_data_a = 16'b1110110010100000;
            14'h5aea: o_data_a = 16'b1110001100001000;
            14'h5aeb: o_data_a = 16'b0000000000000010;
            14'h5aec: o_data_a = 16'b1110110000010000;
            14'h5aed: o_data_a = 16'b0000000000001101;
            14'h5aee: o_data_a = 16'b1110001100001000;
            14'h5aef: o_data_a = 16'b0010000011010110;
            14'h5af0: o_data_a = 16'b1110110000010000;
            14'h5af1: o_data_a = 16'b0000000000001110;
            14'h5af2: o_data_a = 16'b1110001100001000;
            14'h5af3: o_data_a = 16'b0101101011110111;
            14'h5af4: o_data_a = 16'b1110110000010000;
            14'h5af5: o_data_a = 16'b0000000001011111;
            14'h5af6: o_data_a = 16'b1110101010000111;
            14'h5af7: o_data_a = 16'b0000000000000001;
            14'h5af8: o_data_a = 16'b1111110000010000;
            14'h5af9: o_data_a = 16'b0000000000000111;
            14'h5afa: o_data_a = 16'b1110000010010000;
            14'h5afb: o_data_a = 16'b0000000000001101;
            14'h5afc: o_data_a = 16'b1110001100001000;
            14'h5afd: o_data_a = 16'b0000000000000000;
            14'h5afe: o_data_a = 16'b1111110010101000;
            14'h5aff: o_data_a = 16'b1111110000010000;
            14'h5b00: o_data_a = 16'b0000000000001101;
            14'h5b01: o_data_a = 16'b1111110000100000;
            14'h5b02: o_data_a = 16'b1110001100001000;
            14'h5b03: o_data_a = 16'b0000000000000010;
            14'h5b04: o_data_a = 16'b1111110111100000;
            14'h5b05: o_data_a = 16'b1111110000010000;
            14'h5b06: o_data_a = 16'b0000000000000000;
            14'h5b07: o_data_a = 16'b1111110111101000;
            14'h5b08: o_data_a = 16'b1110110010100000;
            14'h5b09: o_data_a = 16'b1110001100001000;
            14'h5b0a: o_data_a = 16'b0000000000000010;
            14'h5b0b: o_data_a = 16'b1111110111100000;
            14'h5b0c: o_data_a = 16'b1110110111100000;
            14'h5b0d: o_data_a = 16'b1111110000010000;
            14'h5b0e: o_data_a = 16'b0000000000000000;
            14'h5b0f: o_data_a = 16'b1111110111101000;
            14'h5b10: o_data_a = 16'b1110110010100000;
            14'h5b11: o_data_a = 16'b1110001100001000;
            14'h5b12: o_data_a = 16'b0000000000000010;
            14'h5b13: o_data_a = 16'b1110110000010000;
            14'h5b14: o_data_a = 16'b0000000000001101;
            14'h5b15: o_data_a = 16'b1110001100001000;
            14'h5b16: o_data_a = 16'b0010000010100111;
            14'h5b17: o_data_a = 16'b1110110000010000;
            14'h5b18: o_data_a = 16'b0000000000001110;
            14'h5b19: o_data_a = 16'b1110001100001000;
            14'h5b1a: o_data_a = 16'b0101101100011110;
            14'h5b1b: o_data_a = 16'b1110110000010000;
            14'h5b1c: o_data_a = 16'b0000000001011111;
            14'h5b1d: o_data_a = 16'b1110101010000111;
            14'h5b1e: o_data_a = 16'b0000000000000001;
            14'h5b1f: o_data_a = 16'b1111110000010000;
            14'h5b20: o_data_a = 16'b0000000000001000;
            14'h5b21: o_data_a = 16'b1110000010010000;
            14'h5b22: o_data_a = 16'b0000000000001101;
            14'h5b23: o_data_a = 16'b1110001100001000;
            14'h5b24: o_data_a = 16'b0000000000000000;
            14'h5b25: o_data_a = 16'b1111110010101000;
            14'h5b26: o_data_a = 16'b1111110000010000;
            14'h5b27: o_data_a = 16'b0000000000001101;
            14'h5b28: o_data_a = 16'b1111110000100000;
            14'h5b29: o_data_a = 16'b1110001100001000;
            14'h5b2a: o_data_a = 16'b0000000000000010;
            14'h5b2b: o_data_a = 16'b1111110000100000;
            14'h5b2c: o_data_a = 16'b1111110000010000;
            14'h5b2d: o_data_a = 16'b0000000000000000;
            14'h5b2e: o_data_a = 16'b1111110111101000;
            14'h5b2f: o_data_a = 16'b1110110010100000;
            14'h5b30: o_data_a = 16'b1110001100001000;
            14'h5b31: o_data_a = 16'b0000000000000000;
            14'h5b32: o_data_a = 16'b1111110111001000;
            14'h5b33: o_data_a = 16'b1111110010100000;
            14'h5b34: o_data_a = 16'b1110111111001000;
            14'h5b35: o_data_a = 16'b0000000000000000;
            14'h5b36: o_data_a = 16'b1111110010100000;
            14'h5b37: o_data_a = 16'b1111110001010000;
            14'h5b38: o_data_a = 16'b1110011111001000;
            14'h5b39: o_data_a = 16'b0101101100111101;
            14'h5b3a: o_data_a = 16'b1110110000010000;
            14'h5b3b: o_data_a = 16'b0000000000010110;
            14'h5b3c: o_data_a = 16'b1110101010000111;
            14'h5b3d: o_data_a = 16'b0000000000000010;
            14'h5b3e: o_data_a = 16'b1111110000100000;
            14'h5b3f: o_data_a = 16'b1111110000010000;
            14'h5b40: o_data_a = 16'b0000000000000000;
            14'h5b41: o_data_a = 16'b1111110111101000;
            14'h5b42: o_data_a = 16'b1110110010100000;
            14'h5b43: o_data_a = 16'b1110001100001000;
            14'h5b44: o_data_a = 16'b0000000100000000;
            14'h5b45: o_data_a = 16'b1110110000010000;
            14'h5b46: o_data_a = 16'b0000000000000000;
            14'h5b47: o_data_a = 16'b1111110111101000;
            14'h5b48: o_data_a = 16'b1110110010100000;
            14'h5b49: o_data_a = 16'b1110001100001000;
            14'h5b4a: o_data_a = 16'b0101101101001110;
            14'h5b4b: o_data_a = 16'b1110110000010000;
            14'h5b4c: o_data_a = 16'b0000000000100110;
            14'h5b4d: o_data_a = 16'b1110101010000111;
            14'h5b4e: o_data_a = 16'b0000000000000000;
            14'h5b4f: o_data_a = 16'b1111110010101000;
            14'h5b50: o_data_a = 16'b1111110000010000;
            14'h5b51: o_data_a = 16'b1110110010100000;
            14'h5b52: o_data_a = 16'b1111000000001000;
            14'h5b53: o_data_a = 16'b0000000000000001;
            14'h5b54: o_data_a = 16'b1111110000010000;
            14'h5b55: o_data_a = 16'b0000000000000111;
            14'h5b56: o_data_a = 16'b1110000010100000;
            14'h5b57: o_data_a = 16'b1111110000010000;
            14'h5b58: o_data_a = 16'b0000000000000000;
            14'h5b59: o_data_a = 16'b1111110111101000;
            14'h5b5a: o_data_a = 16'b1110110010100000;
            14'h5b5b: o_data_a = 16'b1110001100001000;
            14'h5b5c: o_data_a = 16'b0000001000000000;
            14'h5b5d: o_data_a = 16'b1110110000010000;
            14'h5b5e: o_data_a = 16'b0000000000000000;
            14'h5b5f: o_data_a = 16'b1111110111101000;
            14'h5b60: o_data_a = 16'b1110110010100000;
            14'h5b61: o_data_a = 16'b1110001100001000;
            14'h5b62: o_data_a = 16'b0101101101100110;
            14'h5b63: o_data_a = 16'b1110110000010000;
            14'h5b64: o_data_a = 16'b0000000000100110;
            14'h5b65: o_data_a = 16'b1110101010000111;
            14'h5b66: o_data_a = 16'b0000000000000000;
            14'h5b67: o_data_a = 16'b1111110010101000;
            14'h5b68: o_data_a = 16'b1111110000010000;
            14'h5b69: o_data_a = 16'b1110110010100000;
            14'h5b6a: o_data_a = 16'b1111000000001000;
            14'h5b6b: o_data_a = 16'b0000000000000001;
            14'h5b6c: o_data_a = 16'b1111110000010000;
            14'h5b6d: o_data_a = 16'b0000000000001000;
            14'h5b6e: o_data_a = 16'b1110000010100000;
            14'h5b6f: o_data_a = 16'b1111110000010000;
            14'h5b70: o_data_a = 16'b0000000000000000;
            14'h5b71: o_data_a = 16'b1111110111101000;
            14'h5b72: o_data_a = 16'b1110110010100000;
            14'h5b73: o_data_a = 16'b1110001100001000;
            14'h5b74: o_data_a = 16'b0000000000000000;
            14'h5b75: o_data_a = 16'b1111110111001000;
            14'h5b76: o_data_a = 16'b1111110010100000;
            14'h5b77: o_data_a = 16'b1110111111001000;
            14'h5b78: o_data_a = 16'b0000000000000000;
            14'h5b79: o_data_a = 16'b1111110010100000;
            14'h5b7a: o_data_a = 16'b1111110001010000;
            14'h5b7b: o_data_a = 16'b1110011111001000;
            14'h5b7c: o_data_a = 16'b0101101110000000;
            14'h5b7d: o_data_a = 16'b1110110000010000;
            14'h5b7e: o_data_a = 16'b0000000000010110;
            14'h5b7f: o_data_a = 16'b1110101010000111;
            14'h5b80: o_data_a = 16'b0000000000000000;
            14'h5b81: o_data_a = 16'b1111110010101000;
            14'h5b82: o_data_a = 16'b1111110000010000;
            14'h5b83: o_data_a = 16'b1110110010100000;
            14'h5b84: o_data_a = 16'b1111000000001000;
            14'h5b85: o_data_a = 16'b0000000000000000;
            14'h5b86: o_data_a = 16'b1111110010101000;
            14'h5b87: o_data_a = 16'b1111110000010000;
            14'h5b88: o_data_a = 16'b0101101110001100;
            14'h5b89: o_data_a = 16'b1110001100000101;
            14'h5b8a: o_data_a = 16'b0101111001010001;
            14'h5b8b: o_data_a = 16'b1110101010000111;
            14'h5b8c: o_data_a = 16'b0000000000000001;
            14'h5b8d: o_data_a = 16'b1111110000010000;
            14'h5b8e: o_data_a = 16'b0000000000000111;
            14'h5b8f: o_data_a = 16'b1110000010100000;
            14'h5b90: o_data_a = 16'b1111110000010000;
            14'h5b91: o_data_a = 16'b0000000000000000;
            14'h5b92: o_data_a = 16'b1111110111101000;
            14'h5b93: o_data_a = 16'b1110110010100000;
            14'h5b94: o_data_a = 16'b1110001100001000;
            14'h5b95: o_data_a = 16'b0000000000000000;
            14'h5b96: o_data_a = 16'b1111110111001000;
            14'h5b97: o_data_a = 16'b1111110010100000;
            14'h5b98: o_data_a = 16'b1110101010001000;
            14'h5b99: o_data_a = 16'b0000000000000010;
            14'h5b9a: o_data_a = 16'b1110110000010000;
            14'h5b9b: o_data_a = 16'b0000000000001101;
            14'h5b9c: o_data_a = 16'b1110001100001000;
            14'h5b9d: o_data_a = 16'b0010000010100111;
            14'h5b9e: o_data_a = 16'b1110110000010000;
            14'h5b9f: o_data_a = 16'b0000000000001110;
            14'h5ba0: o_data_a = 16'b1110001100001000;
            14'h5ba1: o_data_a = 16'b0101101110100101;
            14'h5ba2: o_data_a = 16'b1110110000010000;
            14'h5ba3: o_data_a = 16'b0000000001011111;
            14'h5ba4: o_data_a = 16'b1110101010000111;
            14'h5ba5: o_data_a = 16'b0000000000000001;
            14'h5ba6: o_data_a = 16'b1111110000010000;
            14'h5ba7: o_data_a = 16'b0000000000000111;
            14'h5ba8: o_data_a = 16'b1110000010010000;
            14'h5ba9: o_data_a = 16'b0000000000001101;
            14'h5baa: o_data_a = 16'b1110001100001000;
            14'h5bab: o_data_a = 16'b0000000000000000;
            14'h5bac: o_data_a = 16'b1111110010101000;
            14'h5bad: o_data_a = 16'b1111110000010000;
            14'h5bae: o_data_a = 16'b0000000000001101;
            14'h5baf: o_data_a = 16'b1111110000100000;
            14'h5bb0: o_data_a = 16'b1110001100001000;
            14'h5bb1: o_data_a = 16'b0000000000000001;
            14'h5bb2: o_data_a = 16'b1111110000010000;
            14'h5bb3: o_data_a = 16'b0000000000001000;
            14'h5bb4: o_data_a = 16'b1110000010100000;
            14'h5bb5: o_data_a = 16'b1111110000010000;
            14'h5bb6: o_data_a = 16'b0000000000000000;
            14'h5bb7: o_data_a = 16'b1111110111101000;
            14'h5bb8: o_data_a = 16'b1110110010100000;
            14'h5bb9: o_data_a = 16'b1110001100001000;
            14'h5bba: o_data_a = 16'b0000000111111111;
            14'h5bbb: o_data_a = 16'b1110110000010000;
            14'h5bbc: o_data_a = 16'b0000000000000000;
            14'h5bbd: o_data_a = 16'b1111110111101000;
            14'h5bbe: o_data_a = 16'b1110110010100000;
            14'h5bbf: o_data_a = 16'b1110001100001000;
            14'h5bc0: o_data_a = 16'b0000000000000010;
            14'h5bc1: o_data_a = 16'b1110110000010000;
            14'h5bc2: o_data_a = 16'b0000000000001101;
            14'h5bc3: o_data_a = 16'b1110001100001000;
            14'h5bc4: o_data_a = 16'b0010000011010110;
            14'h5bc5: o_data_a = 16'b1110110000010000;
            14'h5bc6: o_data_a = 16'b0000000000001110;
            14'h5bc7: o_data_a = 16'b1110001100001000;
            14'h5bc8: o_data_a = 16'b0101101111001100;
            14'h5bc9: o_data_a = 16'b1110110000010000;
            14'h5bca: o_data_a = 16'b0000000001011111;
            14'h5bcb: o_data_a = 16'b1110101010000111;
            14'h5bcc: o_data_a = 16'b0000000000000001;
            14'h5bcd: o_data_a = 16'b1111110000010000;
            14'h5bce: o_data_a = 16'b0000000000001000;
            14'h5bcf: o_data_a = 16'b1110000010010000;
            14'h5bd0: o_data_a = 16'b0000000000001101;
            14'h5bd1: o_data_a = 16'b1110001100001000;
            14'h5bd2: o_data_a = 16'b0000000000000000;
            14'h5bd3: o_data_a = 16'b1111110010101000;
            14'h5bd4: o_data_a = 16'b1111110000010000;
            14'h5bd5: o_data_a = 16'b0000000000001101;
            14'h5bd6: o_data_a = 16'b1111110000100000;
            14'h5bd7: o_data_a = 16'b1110001100001000;
            14'h5bd8: o_data_a = 16'b0000000000000001;
            14'h5bd9: o_data_a = 16'b1111110000010000;
            14'h5bda: o_data_a = 16'b0000000000000111;
            14'h5bdb: o_data_a = 16'b1110000010100000;
            14'h5bdc: o_data_a = 16'b1111110000010000;
            14'h5bdd: o_data_a = 16'b0000000000000000;
            14'h5bde: o_data_a = 16'b1111110111101000;
            14'h5bdf: o_data_a = 16'b1110110010100000;
            14'h5be0: o_data_a = 16'b1110001100001000;
            14'h5be1: o_data_a = 16'b0000000000010000;
            14'h5be2: o_data_a = 16'b1110110000010000;
            14'h5be3: o_data_a = 16'b0000000000000000;
            14'h5be4: o_data_a = 16'b1111110111101000;
            14'h5be5: o_data_a = 16'b1110110010100000;
            14'h5be6: o_data_a = 16'b1110001100001000;
            14'h5be7: o_data_a = 16'b0000000000000010;
            14'h5be8: o_data_a = 16'b1110110000010000;
            14'h5be9: o_data_a = 16'b0000000000001101;
            14'h5bea: o_data_a = 16'b1110001100001000;
            14'h5beb: o_data_a = 16'b0001110001110111;
            14'h5bec: o_data_a = 16'b1110110000010000;
            14'h5bed: o_data_a = 16'b0000000000001110;
            14'h5bee: o_data_a = 16'b1110001100001000;
            14'h5bef: o_data_a = 16'b0101101111110011;
            14'h5bf0: o_data_a = 16'b1110110000010000;
            14'h5bf1: o_data_a = 16'b0000000001011111;
            14'h5bf2: o_data_a = 16'b1110101010000111;
            14'h5bf3: o_data_a = 16'b0000000000000000;
            14'h5bf4: o_data_a = 16'b1111110010101000;
            14'h5bf5: o_data_a = 16'b1111110000010000;
            14'h5bf6: o_data_a = 16'b0000000000000001;
            14'h5bf7: o_data_a = 16'b1111110111100000;
            14'h5bf8: o_data_a = 16'b1110001100001000;
            14'h5bf9: o_data_a = 16'b0000000000000001;
            14'h5bfa: o_data_a = 16'b1111110000010000;
            14'h5bfb: o_data_a = 16'b0000000000000111;
            14'h5bfc: o_data_a = 16'b1110000010100000;
            14'h5bfd: o_data_a = 16'b1111110000010000;
            14'h5bfe: o_data_a = 16'b0000000000000000;
            14'h5bff: o_data_a = 16'b1111110111101000;
            14'h5c00: o_data_a = 16'b1110110010100000;
            14'h5c01: o_data_a = 16'b1110001100001000;
            14'h5c02: o_data_a = 16'b0000000000000001;
            14'h5c03: o_data_a = 16'b1111110111100000;
            14'h5c04: o_data_a = 16'b1111110000010000;
            14'h5c05: o_data_a = 16'b0000000000000000;
            14'h5c06: o_data_a = 16'b1111110111101000;
            14'h5c07: o_data_a = 16'b1110110010100000;
            14'h5c08: o_data_a = 16'b1110001100001000;
            14'h5c09: o_data_a = 16'b0000000000010000;
            14'h5c0a: o_data_a = 16'b1110110000010000;
            14'h5c0b: o_data_a = 16'b0000000000000000;
            14'h5c0c: o_data_a = 16'b1111110111101000;
            14'h5c0d: o_data_a = 16'b1110110010100000;
            14'h5c0e: o_data_a = 16'b1110001100001000;
            14'h5c0f: o_data_a = 16'b0000000000000010;
            14'h5c10: o_data_a = 16'b1110110000010000;
            14'h5c11: o_data_a = 16'b0000000000001101;
            14'h5c12: o_data_a = 16'b1110001100001000;
            14'h5c13: o_data_a = 16'b0001101010100110;
            14'h5c14: o_data_a = 16'b1110110000010000;
            14'h5c15: o_data_a = 16'b0000000000001110;
            14'h5c16: o_data_a = 16'b1110001100001000;
            14'h5c17: o_data_a = 16'b0101110000011011;
            14'h5c18: o_data_a = 16'b1110110000010000;
            14'h5c19: o_data_a = 16'b0000000001011111;
            14'h5c1a: o_data_a = 16'b1110101010000111;
            14'h5c1b: o_data_a = 16'b0000000000000000;
            14'h5c1c: o_data_a = 16'b1111110010101000;
            14'h5c1d: o_data_a = 16'b1111110000010000;
            14'h5c1e: o_data_a = 16'b1110110010100000;
            14'h5c1f: o_data_a = 16'b1111000111001000;
            14'h5c20: o_data_a = 16'b0000000000000001;
            14'h5c21: o_data_a = 16'b1111110000010000;
            14'h5c22: o_data_a = 16'b0000000000001001;
            14'h5c23: o_data_a = 16'b1110000010010000;
            14'h5c24: o_data_a = 16'b0000000000001101;
            14'h5c25: o_data_a = 16'b1110001100001000;
            14'h5c26: o_data_a = 16'b0000000000000000;
            14'h5c27: o_data_a = 16'b1111110010101000;
            14'h5c28: o_data_a = 16'b1111110000010000;
            14'h5c29: o_data_a = 16'b0000000000001101;
            14'h5c2a: o_data_a = 16'b1111110000100000;
            14'h5c2b: o_data_a = 16'b1110001100001000;
            14'h5c2c: o_data_a = 16'b0000000000000001;
            14'h5c2d: o_data_a = 16'b1111110000010000;
            14'h5c2e: o_data_a = 16'b0000000000001000;
            14'h5c2f: o_data_a = 16'b1110000010100000;
            14'h5c30: o_data_a = 16'b1111110000010000;
            14'h5c31: o_data_a = 16'b0000000000000000;
            14'h5c32: o_data_a = 16'b1111110111101000;
            14'h5c33: o_data_a = 16'b1110110010100000;
            14'h5c34: o_data_a = 16'b1110001100001000;
            14'h5c35: o_data_a = 16'b0000000000010000;
            14'h5c36: o_data_a = 16'b1110110000010000;
            14'h5c37: o_data_a = 16'b0000000000000000;
            14'h5c38: o_data_a = 16'b1111110111101000;
            14'h5c39: o_data_a = 16'b1110110010100000;
            14'h5c3a: o_data_a = 16'b1110001100001000;
            14'h5c3b: o_data_a = 16'b0000000000000010;
            14'h5c3c: o_data_a = 16'b1110110000010000;
            14'h5c3d: o_data_a = 16'b0000000000001101;
            14'h5c3e: o_data_a = 16'b1110001100001000;
            14'h5c3f: o_data_a = 16'b0001110001110111;
            14'h5c40: o_data_a = 16'b1110110000010000;
            14'h5c41: o_data_a = 16'b0000000000001110;
            14'h5c42: o_data_a = 16'b1110001100001000;
            14'h5c43: o_data_a = 16'b0101110001000111;
            14'h5c44: o_data_a = 16'b1110110000010000;
            14'h5c45: o_data_a = 16'b0000000001011111;
            14'h5c46: o_data_a = 16'b1110101010000111;
            14'h5c47: o_data_a = 16'b0000000000000000;
            14'h5c48: o_data_a = 16'b1111110010101000;
            14'h5c49: o_data_a = 16'b1111110000010000;
            14'h5c4a: o_data_a = 16'b0000000000000001;
            14'h5c4b: o_data_a = 16'b1111110111100000;
            14'h5c4c: o_data_a = 16'b1110110111100000;
            14'h5c4d: o_data_a = 16'b1110001100001000;
            14'h5c4e: o_data_a = 16'b0000000000000001;
            14'h5c4f: o_data_a = 16'b1111110000010000;
            14'h5c50: o_data_a = 16'b0000000000001000;
            14'h5c51: o_data_a = 16'b1110000010100000;
            14'h5c52: o_data_a = 16'b1111110000010000;
            14'h5c53: o_data_a = 16'b0000000000000000;
            14'h5c54: o_data_a = 16'b1111110111101000;
            14'h5c55: o_data_a = 16'b1110110010100000;
            14'h5c56: o_data_a = 16'b1110001100001000;
            14'h5c57: o_data_a = 16'b0000000000000001;
            14'h5c58: o_data_a = 16'b1111110111100000;
            14'h5c59: o_data_a = 16'b1110110111100000;
            14'h5c5a: o_data_a = 16'b1111110000010000;
            14'h5c5b: o_data_a = 16'b0000000000000000;
            14'h5c5c: o_data_a = 16'b1111110111101000;
            14'h5c5d: o_data_a = 16'b1110110010100000;
            14'h5c5e: o_data_a = 16'b1110001100001000;
            14'h5c5f: o_data_a = 16'b0000000000010000;
            14'h5c60: o_data_a = 16'b1110110000010000;
            14'h5c61: o_data_a = 16'b0000000000000000;
            14'h5c62: o_data_a = 16'b1111110111101000;
            14'h5c63: o_data_a = 16'b1110110010100000;
            14'h5c64: o_data_a = 16'b1110001100001000;
            14'h5c65: o_data_a = 16'b0000000000000010;
            14'h5c66: o_data_a = 16'b1110110000010000;
            14'h5c67: o_data_a = 16'b0000000000001101;
            14'h5c68: o_data_a = 16'b1110001100001000;
            14'h5c69: o_data_a = 16'b0001101010100110;
            14'h5c6a: o_data_a = 16'b1110110000010000;
            14'h5c6b: o_data_a = 16'b0000000000001110;
            14'h5c6c: o_data_a = 16'b1110001100001000;
            14'h5c6d: o_data_a = 16'b0101110001110001;
            14'h5c6e: o_data_a = 16'b1110110000010000;
            14'h5c6f: o_data_a = 16'b0000000001011111;
            14'h5c70: o_data_a = 16'b1110101010000111;
            14'h5c71: o_data_a = 16'b0000000000000000;
            14'h5c72: o_data_a = 16'b1111110010101000;
            14'h5c73: o_data_a = 16'b1111110000010000;
            14'h5c74: o_data_a = 16'b1110110010100000;
            14'h5c75: o_data_a = 16'b1111000111001000;
            14'h5c76: o_data_a = 16'b0000000000000001;
            14'h5c77: o_data_a = 16'b1111110000010000;
            14'h5c78: o_data_a = 16'b0000000000001010;
            14'h5c79: o_data_a = 16'b1110000010010000;
            14'h5c7a: o_data_a = 16'b0000000000001101;
            14'h5c7b: o_data_a = 16'b1110001100001000;
            14'h5c7c: o_data_a = 16'b0000000000000000;
            14'h5c7d: o_data_a = 16'b1111110010101000;
            14'h5c7e: o_data_a = 16'b1111110000010000;
            14'h5c7f: o_data_a = 16'b0000000000001101;
            14'h5c80: o_data_a = 16'b1111110000100000;
            14'h5c81: o_data_a = 16'b1110001100001000;
            14'h5c82: o_data_a = 16'b0000000000000001;
            14'h5c83: o_data_a = 16'b1111110000010000;
            14'h5c84: o_data_a = 16'b0000000000001001;
            14'h5c85: o_data_a = 16'b1110000010100000;
            14'h5c86: o_data_a = 16'b1111110000010000;
            14'h5c87: o_data_a = 16'b0000000000000000;
            14'h5c88: o_data_a = 16'b1111110111101000;
            14'h5c89: o_data_a = 16'b1110110010100000;
            14'h5c8a: o_data_a = 16'b1110001100001000;
            14'h5c8b: o_data_a = 16'b0000000000011101;
            14'h5c8c: o_data_a = 16'b1111110000010000;
            14'h5c8d: o_data_a = 16'b0000000000000000;
            14'h5c8e: o_data_a = 16'b1111110111101000;
            14'h5c8f: o_data_a = 16'b1110110010100000;
            14'h5c90: o_data_a = 16'b1110001100001000;
            14'h5c91: o_data_a = 16'b0000000000000000;
            14'h5c92: o_data_a = 16'b1111110010101000;
            14'h5c93: o_data_a = 16'b1111110000010000;
            14'h5c94: o_data_a = 16'b1110110010100000;
            14'h5c95: o_data_a = 16'b1111000010001000;
            14'h5c96: o_data_a = 16'b0000000000000000;
            14'h5c97: o_data_a = 16'b1111110010101000;
            14'h5c98: o_data_a = 16'b1111110000010000;
            14'h5c99: o_data_a = 16'b0000000000000100;
            14'h5c9a: o_data_a = 16'b1110001100001000;
            14'h5c9b: o_data_a = 16'b0000000000000100;
            14'h5c9c: o_data_a = 16'b1111110000100000;
            14'h5c9d: o_data_a = 16'b1111110000010000;
            14'h5c9e: o_data_a = 16'b0000000000000000;
            14'h5c9f: o_data_a = 16'b1111110111101000;
            14'h5ca0: o_data_a = 16'b1110110010100000;
            14'h5ca1: o_data_a = 16'b1110001100001000;
            14'h5ca2: o_data_a = 16'b0000000000000000;
            14'h5ca3: o_data_a = 16'b1111110111001000;
            14'h5ca4: o_data_a = 16'b1111110010100000;
            14'h5ca5: o_data_a = 16'b1110111111001000;
            14'h5ca6: o_data_a = 16'b0000000000000000;
            14'h5ca7: o_data_a = 16'b1111110010101000;
            14'h5ca8: o_data_a = 16'b1111110000010000;
            14'h5ca9: o_data_a = 16'b1110110010100000;
            14'h5caa: o_data_a = 16'b1111000111001000;
            14'h5cab: o_data_a = 16'b0000000000000000;
            14'h5cac: o_data_a = 16'b1111110010100000;
            14'h5cad: o_data_a = 16'b1111110001001000;
            14'h5cae: o_data_a = 16'b0000000000000000;
            14'h5caf: o_data_a = 16'b1111110010101000;
            14'h5cb0: o_data_a = 16'b1111110000010000;
            14'h5cb1: o_data_a = 16'b0000000000000001;
            14'h5cb2: o_data_a = 16'b1111110111100000;
            14'h5cb3: o_data_a = 16'b1110110111100000;
            14'h5cb4: o_data_a = 16'b1110110111100000;
            14'h5cb5: o_data_a = 16'b1110110111100000;
            14'h5cb6: o_data_a = 16'b1110110111100000;
            14'h5cb7: o_data_a = 16'b1110001100001000;
            14'h5cb8: o_data_a = 16'b0000000000000001;
            14'h5cb9: o_data_a = 16'b1111110000010000;
            14'h5cba: o_data_a = 16'b0000000000001010;
            14'h5cbb: o_data_a = 16'b1110000010100000;
            14'h5cbc: o_data_a = 16'b1111110000010000;
            14'h5cbd: o_data_a = 16'b0000000000000000;
            14'h5cbe: o_data_a = 16'b1111110111101000;
            14'h5cbf: o_data_a = 16'b1110110010100000;
            14'h5cc0: o_data_a = 16'b1110001100001000;
            14'h5cc1: o_data_a = 16'b0000000000000000;
            14'h5cc2: o_data_a = 16'b1111110111001000;
            14'h5cc3: o_data_a = 16'b1111110010100000;
            14'h5cc4: o_data_a = 16'b1110111111001000;
            14'h5cc5: o_data_a = 16'b0000000000000000;
            14'h5cc6: o_data_a = 16'b1111110010101000;
            14'h5cc7: o_data_a = 16'b1111110000010000;
            14'h5cc8: o_data_a = 16'b1110110010100000;
            14'h5cc9: o_data_a = 16'b1111000010001000;
            14'h5cca: o_data_a = 16'b0000000000011101;
            14'h5ccb: o_data_a = 16'b1111110000010000;
            14'h5ccc: o_data_a = 16'b0000000000000000;
            14'h5ccd: o_data_a = 16'b1111110111101000;
            14'h5cce: o_data_a = 16'b1110110010100000;
            14'h5ccf: o_data_a = 16'b1110001100001000;
            14'h5cd0: o_data_a = 16'b0000000000000000;
            14'h5cd1: o_data_a = 16'b1111110010101000;
            14'h5cd2: o_data_a = 16'b1111110000010000;
            14'h5cd3: o_data_a = 16'b1110110010100000;
            14'h5cd4: o_data_a = 16'b1111000010001000;
            14'h5cd5: o_data_a = 16'b0000000000000000;
            14'h5cd6: o_data_a = 16'b1111110010101000;
            14'h5cd7: o_data_a = 16'b1111110000010000;
            14'h5cd8: o_data_a = 16'b0000000000000100;
            14'h5cd9: o_data_a = 16'b1110001100001000;
            14'h5cda: o_data_a = 16'b0000000000000100;
            14'h5cdb: o_data_a = 16'b1111110000100000;
            14'h5cdc: o_data_a = 16'b1111110000010000;
            14'h5cdd: o_data_a = 16'b0000000000000000;
            14'h5cde: o_data_a = 16'b1111110111101000;
            14'h5cdf: o_data_a = 16'b1110110010100000;
            14'h5ce0: o_data_a = 16'b1110001100001000;
            14'h5ce1: o_data_a = 16'b0000000000000000;
            14'h5ce2: o_data_a = 16'b1111110111001000;
            14'h5ce3: o_data_a = 16'b1111110010100000;
            14'h5ce4: o_data_a = 16'b1110111111001000;
            14'h5ce5: o_data_a = 16'b0000000000000000;
            14'h5ce6: o_data_a = 16'b1111110010101000;
            14'h5ce7: o_data_a = 16'b1111110000010000;
            14'h5ce8: o_data_a = 16'b1110110010100000;
            14'h5ce9: o_data_a = 16'b1111000111001000;
            14'h5cea: o_data_a = 16'b0000000000000000;
            14'h5ceb: o_data_a = 16'b1111110010101000;
            14'h5cec: o_data_a = 16'b1111110000010000;
            14'h5ced: o_data_a = 16'b0000000000000001;
            14'h5cee: o_data_a = 16'b1111110111100000;
            14'h5cef: o_data_a = 16'b1110110111100000;
            14'h5cf0: o_data_a = 16'b1110110111100000;
            14'h5cf1: o_data_a = 16'b1110110111100000;
            14'h5cf2: o_data_a = 16'b1110001100001000;
            14'h5cf3: o_data_a = 16'b0000000000000010;
            14'h5cf4: o_data_a = 16'b1111110000100000;
            14'h5cf5: o_data_a = 16'b1111110000010000;
            14'h5cf6: o_data_a = 16'b0000000000000000;
            14'h5cf7: o_data_a = 16'b1111110111101000;
            14'h5cf8: o_data_a = 16'b1110110010100000;
            14'h5cf9: o_data_a = 16'b1110001100001000;
            14'h5cfa: o_data_a = 16'b0000000000100000;
            14'h5cfb: o_data_a = 16'b1110110000010000;
            14'h5cfc: o_data_a = 16'b0000000000000000;
            14'h5cfd: o_data_a = 16'b1111110111101000;
            14'h5cfe: o_data_a = 16'b1110110010100000;
            14'h5cff: o_data_a = 16'b1110001100001000;
            14'h5d00: o_data_a = 16'b0000000000000010;
            14'h5d01: o_data_a = 16'b1110110000010000;
            14'h5d02: o_data_a = 16'b0000000000001101;
            14'h5d03: o_data_a = 16'b1110001100001000;
            14'h5d04: o_data_a = 16'b0001101010100110;
            14'h5d05: o_data_a = 16'b1110110000010000;
            14'h5d06: o_data_a = 16'b0000000000001110;
            14'h5d07: o_data_a = 16'b1110001100001000;
            14'h5d08: o_data_a = 16'b0101110100001100;
            14'h5d09: o_data_a = 16'b1110110000010000;
            14'h5d0a: o_data_a = 16'b0000000001011111;
            14'h5d0b: o_data_a = 16'b1110101010000111;
            14'h5d0c: o_data_a = 16'b0000000000000001;
            14'h5d0d: o_data_a = 16'b1111110111100000;
            14'h5d0e: o_data_a = 16'b1111110000010000;
            14'h5d0f: o_data_a = 16'b0000000000000000;
            14'h5d10: o_data_a = 16'b1111110111101000;
            14'h5d11: o_data_a = 16'b1110110010100000;
            14'h5d12: o_data_a = 16'b1110001100001000;
            14'h5d13: o_data_a = 16'b0000000000000000;
            14'h5d14: o_data_a = 16'b1111110010101000;
            14'h5d15: o_data_a = 16'b1111110000010000;
            14'h5d16: o_data_a = 16'b1110110010100000;
            14'h5d17: o_data_a = 16'b1111000010001000;
            14'h5d18: o_data_a = 16'b0000000000000000;
            14'h5d19: o_data_a = 16'b1111110010101000;
            14'h5d1a: o_data_a = 16'b1111110000010000;
            14'h5d1b: o_data_a = 16'b0000000000000001;
            14'h5d1c: o_data_a = 16'b1111110000100000;
            14'h5d1d: o_data_a = 16'b1110001100001000;
            14'h5d1e: o_data_a = 16'b0000000000000001;
            14'h5d1f: o_data_a = 16'b1111110111100000;
            14'h5d20: o_data_a = 16'b1110110111100000;
            14'h5d21: o_data_a = 16'b1111110000010000;
            14'h5d22: o_data_a = 16'b0000000000000000;
            14'h5d23: o_data_a = 16'b1111110111101000;
            14'h5d24: o_data_a = 16'b1110110010100000;
            14'h5d25: o_data_a = 16'b1110001100001000;
            14'h5d26: o_data_a = 16'b0000000000000001;
            14'h5d27: o_data_a = 16'b1111110111100000;
            14'h5d28: o_data_a = 16'b1111110000010000;
            14'h5d29: o_data_a = 16'b0000000000000000;
            14'h5d2a: o_data_a = 16'b1111110111101000;
            14'h5d2b: o_data_a = 16'b1110110010100000;
            14'h5d2c: o_data_a = 16'b1110001100001000;
            14'h5d2d: o_data_a = 16'b0000000000000000;
            14'h5d2e: o_data_a = 16'b1111110010101000;
            14'h5d2f: o_data_a = 16'b1111110000010000;
            14'h5d30: o_data_a = 16'b1110110010100000;
            14'h5d31: o_data_a = 16'b1111000111001000;
            14'h5d32: o_data_a = 16'b0000000000000000;
            14'h5d33: o_data_a = 16'b1111110010101000;
            14'h5d34: o_data_a = 16'b1111110000010000;
            14'h5d35: o_data_a = 16'b0000000000000001;
            14'h5d36: o_data_a = 16'b1111110111100000;
            14'h5d37: o_data_a = 16'b1110110111100000;
            14'h5d38: o_data_a = 16'b1110110111100000;
            14'h5d39: o_data_a = 16'b1110110111100000;
            14'h5d3a: o_data_a = 16'b1110110111100000;
            14'h5d3b: o_data_a = 16'b1110110111100000;
            14'h5d3c: o_data_a = 16'b1110001100001000;
            14'h5d3d: o_data_a = 16'b0000000000000001;
            14'h5d3e: o_data_a = 16'b1111110000100000;
            14'h5d3f: o_data_a = 16'b1111110000010000;
            14'h5d40: o_data_a = 16'b0000000000000000;
            14'h5d41: o_data_a = 16'b1111110111101000;
            14'h5d42: o_data_a = 16'b1110110010100000;
            14'h5d43: o_data_a = 16'b1110001100001000;
            14'h5d44: o_data_a = 16'b0000000000000001;
            14'h5d45: o_data_a = 16'b1111110000010000;
            14'h5d46: o_data_a = 16'b0000000000000110;
            14'h5d47: o_data_a = 16'b1110000010100000;
            14'h5d48: o_data_a = 16'b1111110000010000;
            14'h5d49: o_data_a = 16'b0000000000000000;
            14'h5d4a: o_data_a = 16'b1111110111101000;
            14'h5d4b: o_data_a = 16'b1110110010100000;
            14'h5d4c: o_data_a = 16'b1110001100001000;
            14'h5d4d: o_data_a = 16'b0000000000000000;
            14'h5d4e: o_data_a = 16'b1111110010101000;
            14'h5d4f: o_data_a = 16'b1111110000010000;
            14'h5d50: o_data_a = 16'b1110110010100000;
            14'h5d51: o_data_a = 16'b1111000010001000;
            14'h5d52: o_data_a = 16'b0000000000000000;
            14'h5d53: o_data_a = 16'b1111110010101000;
            14'h5d54: o_data_a = 16'b1111110000010000;
            14'h5d55: o_data_a = 16'b0000000000000001;
            14'h5d56: o_data_a = 16'b1111110111100000;
            14'h5d57: o_data_a = 16'b1110110111100000;
            14'h5d58: o_data_a = 16'b1110110111100000;
            14'h5d59: o_data_a = 16'b1110001100001000;
            14'h5d5a: o_data_a = 16'b0000000000000001;
            14'h5d5b: o_data_a = 16'b1111110000010000;
            14'h5d5c: o_data_a = 16'b0000000000000110;
            14'h5d5d: o_data_a = 16'b1110000010100000;
            14'h5d5e: o_data_a = 16'b1111110000010000;
            14'h5d5f: o_data_a = 16'b0000000000000000;
            14'h5d60: o_data_a = 16'b1111110111101000;
            14'h5d61: o_data_a = 16'b1110110010100000;
            14'h5d62: o_data_a = 16'b1110001100001000;
            14'h5d63: o_data_a = 16'b0000000000000000;
            14'h5d64: o_data_a = 16'b1111110111001000;
            14'h5d65: o_data_a = 16'b1111110010100000;
            14'h5d66: o_data_a = 16'b1110101010001000;
            14'h5d67: o_data_a = 16'b0101110101101011;
            14'h5d68: o_data_a = 16'b1110110000010000;
            14'h5d69: o_data_a = 16'b0000000000000110;
            14'h5d6a: o_data_a = 16'b1110101010000111;
            14'h5d6b: o_data_a = 16'b0000000000000000;
            14'h5d6c: o_data_a = 16'b1111110010101000;
            14'h5d6d: o_data_a = 16'b1111110000010000;
            14'h5d6e: o_data_a = 16'b0101110101110010;
            14'h5d6f: o_data_a = 16'b1110001100000101;
            14'h5d70: o_data_a = 16'b0101110110100011;
            14'h5d71: o_data_a = 16'b1110101010000111;
            14'h5d72: o_data_a = 16'b0000000000000001;
            14'h5d73: o_data_a = 16'b1111110000100000;
            14'h5d74: o_data_a = 16'b1111110000010000;
            14'h5d75: o_data_a = 16'b0000000000000000;
            14'h5d76: o_data_a = 16'b1111110111101000;
            14'h5d77: o_data_a = 16'b1110110010100000;
            14'h5d78: o_data_a = 16'b1110001100001000;
            14'h5d79: o_data_a = 16'b0000000000000001;
            14'h5d7a: o_data_a = 16'b1111110000010000;
            14'h5d7b: o_data_a = 16'b0000000000000100;
            14'h5d7c: o_data_a = 16'b1110000010100000;
            14'h5d7d: o_data_a = 16'b1111110000010000;
            14'h5d7e: o_data_a = 16'b0000000000000000;
            14'h5d7f: o_data_a = 16'b1111110111101000;
            14'h5d80: o_data_a = 16'b1110110010100000;
            14'h5d81: o_data_a = 16'b1110001100001000;
            14'h5d82: o_data_a = 16'b0000000000000001;
            14'h5d83: o_data_a = 16'b1111110000010000;
            14'h5d84: o_data_a = 16'b0000000000000101;
            14'h5d85: o_data_a = 16'b1110000010100000;
            14'h5d86: o_data_a = 16'b1111110000010000;
            14'h5d87: o_data_a = 16'b0000000000000000;
            14'h5d88: o_data_a = 16'b1111110111101000;
            14'h5d89: o_data_a = 16'b1110110010100000;
            14'h5d8a: o_data_a = 16'b1110001100001000;
            14'h5d8b: o_data_a = 16'b0000000000000000;
            14'h5d8c: o_data_a = 16'b1111110010101000;
            14'h5d8d: o_data_a = 16'b1111110000010000;
            14'h5d8e: o_data_a = 16'b1110110010100000;
            14'h5d8f: o_data_a = 16'b1111000000001000;
            14'h5d90: o_data_a = 16'b0000000000000010;
            14'h5d91: o_data_a = 16'b1110110000010000;
            14'h5d92: o_data_a = 16'b0000000000001101;
            14'h5d93: o_data_a = 16'b1110001100001000;
            14'h5d94: o_data_a = 16'b0101000011011101;
            14'h5d95: o_data_a = 16'b1110110000010000;
            14'h5d96: o_data_a = 16'b0000000000001110;
            14'h5d97: o_data_a = 16'b1110001100001000;
            14'h5d98: o_data_a = 16'b0101110110011100;
            14'h5d99: o_data_a = 16'b1110110000010000;
            14'h5d9a: o_data_a = 16'b0000000001011111;
            14'h5d9b: o_data_a = 16'b1110101010000111;
            14'h5d9c: o_data_a = 16'b0000000000000000;
            14'h5d9d: o_data_a = 16'b1111110010101000;
            14'h5d9e: o_data_a = 16'b1111110000010000;
            14'h5d9f: o_data_a = 16'b0000000000000101;
            14'h5da0: o_data_a = 16'b1110001100001000;
            14'h5da1: o_data_a = 16'b0101111001010001;
            14'h5da2: o_data_a = 16'b1110101010000111;
            14'h5da3: o_data_a = 16'b0000000000000001;
            14'h5da4: o_data_a = 16'b1111110000100000;
            14'h5da5: o_data_a = 16'b1111110000010000;
            14'h5da6: o_data_a = 16'b0000000000000000;
            14'h5da7: o_data_a = 16'b1111110111101000;
            14'h5da8: o_data_a = 16'b1110110010100000;
            14'h5da9: o_data_a = 16'b1110001100001000;
            14'h5daa: o_data_a = 16'b0000000000000001;
            14'h5dab: o_data_a = 16'b1111110000010000;
            14'h5dac: o_data_a = 16'b0000000000000101;
            14'h5dad: o_data_a = 16'b1110000010100000;
            14'h5dae: o_data_a = 16'b1111110000010000;
            14'h5daf: o_data_a = 16'b0000000000000000;
            14'h5db0: o_data_a = 16'b1111110111101000;
            14'h5db1: o_data_a = 16'b1110110010100000;
            14'h5db2: o_data_a = 16'b1110001100001000;
            14'h5db3: o_data_a = 16'b0000000000000010;
            14'h5db4: o_data_a = 16'b1110110000010000;
            14'h5db5: o_data_a = 16'b0000000000001101;
            14'h5db6: o_data_a = 16'b1110001100001000;
            14'h5db7: o_data_a = 16'b0101000011011101;
            14'h5db8: o_data_a = 16'b1110110000010000;
            14'h5db9: o_data_a = 16'b0000000000001110;
            14'h5dba: o_data_a = 16'b1110001100001000;
            14'h5dbb: o_data_a = 16'b0101110110111111;
            14'h5dbc: o_data_a = 16'b1110110000010000;
            14'h5dbd: o_data_a = 16'b0000000001011111;
            14'h5dbe: o_data_a = 16'b1110101010000111;
            14'h5dbf: o_data_a = 16'b0000000000000000;
            14'h5dc0: o_data_a = 16'b1111110010101000;
            14'h5dc1: o_data_a = 16'b1111110000010000;
            14'h5dc2: o_data_a = 16'b0000000000000101;
            14'h5dc3: o_data_a = 16'b1110001100001000;
            14'h5dc4: o_data_a = 16'b0000000000000001;
            14'h5dc5: o_data_a = 16'b1111110000100000;
            14'h5dc6: o_data_a = 16'b1111110000010000;
            14'h5dc7: o_data_a = 16'b0000000000000000;
            14'h5dc8: o_data_a = 16'b1111110111101000;
            14'h5dc9: o_data_a = 16'b1110110010100000;
            14'h5dca: o_data_a = 16'b1110001100001000;
            14'h5dcb: o_data_a = 16'b0000000000000000;
            14'h5dcc: o_data_a = 16'b1111110111001000;
            14'h5dcd: o_data_a = 16'b1111110010100000;
            14'h5dce: o_data_a = 16'b1110111111001000;
            14'h5dcf: o_data_a = 16'b0000000000000000;
            14'h5dd0: o_data_a = 16'b1111110010101000;
            14'h5dd1: o_data_a = 16'b1111110000010000;
            14'h5dd2: o_data_a = 16'b1110110010100000;
            14'h5dd3: o_data_a = 16'b1111000010001000;
            14'h5dd4: o_data_a = 16'b0000000000000000;
            14'h5dd5: o_data_a = 16'b1111110010101000;
            14'h5dd6: o_data_a = 16'b1111110000010000;
            14'h5dd7: o_data_a = 16'b0000000000000001;
            14'h5dd8: o_data_a = 16'b1111110000100000;
            14'h5dd9: o_data_a = 16'b1110001100001000;
            14'h5dda: o_data_a = 16'b0000000000000001;
            14'h5ddb: o_data_a = 16'b1111110000100000;
            14'h5ddc: o_data_a = 16'b1111110000010000;
            14'h5ddd: o_data_a = 16'b0000000000000000;
            14'h5dde: o_data_a = 16'b1111110111101000;
            14'h5ddf: o_data_a = 16'b1110110010100000;
            14'h5de0: o_data_a = 16'b1110001100001000;
            14'h5de1: o_data_a = 16'b0000000000000001;
            14'h5de2: o_data_a = 16'b1111110000010000;
            14'h5de3: o_data_a = 16'b0000000000000011;
            14'h5de4: o_data_a = 16'b1110000010100000;
            14'h5de5: o_data_a = 16'b1111110000010000;
            14'h5de6: o_data_a = 16'b0000000000000000;
            14'h5de7: o_data_a = 16'b1111110111101000;
            14'h5de8: o_data_a = 16'b1110110010100000;
            14'h5de9: o_data_a = 16'b1110001100001000;
            14'h5dea: o_data_a = 16'b0101110111101110;
            14'h5deb: o_data_a = 16'b1110110000010000;
            14'h5dec: o_data_a = 16'b0000000000100110;
            14'h5ded: o_data_a = 16'b1110101010000111;
            14'h5dee: o_data_a = 16'b0000000000000000;
            14'h5def: o_data_a = 16'b1111110010100000;
            14'h5df0: o_data_a = 16'b1111110001001000;
            14'h5df1: o_data_a = 16'b0000000000000000;
            14'h5df2: o_data_a = 16'b1111110010101000;
            14'h5df3: o_data_a = 16'b1111110000010000;
            14'h5df4: o_data_a = 16'b0101111000101110;
            14'h5df5: o_data_a = 16'b1110001100000101;
            14'h5df6: o_data_a = 16'b0000000000000001;
            14'h5df7: o_data_a = 16'b1111110000100000;
            14'h5df8: o_data_a = 16'b1111110000010000;
            14'h5df9: o_data_a = 16'b0000000000000000;
            14'h5dfa: o_data_a = 16'b1111110111101000;
            14'h5dfb: o_data_a = 16'b1110110010100000;
            14'h5dfc: o_data_a = 16'b1110001100001000;
            14'h5dfd: o_data_a = 16'b0000000000000000;
            14'h5dfe: o_data_a = 16'b1111110111001000;
            14'h5dff: o_data_a = 16'b1111110010100000;
            14'h5e00: o_data_a = 16'b1110111111001000;
            14'h5e01: o_data_a = 16'b0000000000000000;
            14'h5e02: o_data_a = 16'b1111110010100000;
            14'h5e03: o_data_a = 16'b1111110001010000;
            14'h5e04: o_data_a = 16'b1110011111001000;
            14'h5e05: o_data_a = 16'b0000000000000010;
            14'h5e06: o_data_a = 16'b1110110000010000;
            14'h5e07: o_data_a = 16'b0000000000001101;
            14'h5e08: o_data_a = 16'b1110001100001000;
            14'h5e09: o_data_a = 16'b0101000011011101;
            14'h5e0a: o_data_a = 16'b1110110000010000;
            14'h5e0b: o_data_a = 16'b0000000000001110;
            14'h5e0c: o_data_a = 16'b1110001100001000;
            14'h5e0d: o_data_a = 16'b0101111000010001;
            14'h5e0e: o_data_a = 16'b1110110000010000;
            14'h5e0f: o_data_a = 16'b0000000001011111;
            14'h5e10: o_data_a = 16'b1110101010000111;
            14'h5e11: o_data_a = 16'b0000000000000000;
            14'h5e12: o_data_a = 16'b1111110010101000;
            14'h5e13: o_data_a = 16'b1111110000010000;
            14'h5e14: o_data_a = 16'b0000000000000101;
            14'h5e15: o_data_a = 16'b1110001100001000;
            14'h5e16: o_data_a = 16'b0000000000000001;
            14'h5e17: o_data_a = 16'b1111110000100000;
            14'h5e18: o_data_a = 16'b1111110000010000;
            14'h5e19: o_data_a = 16'b0000000000000000;
            14'h5e1a: o_data_a = 16'b1111110111101000;
            14'h5e1b: o_data_a = 16'b1110110010100000;
            14'h5e1c: o_data_a = 16'b1110001100001000;
            14'h5e1d: o_data_a = 16'b0000000000000000;
            14'h5e1e: o_data_a = 16'b1111110111001000;
            14'h5e1f: o_data_a = 16'b1111110010100000;
            14'h5e20: o_data_a = 16'b1110111111001000;
            14'h5e21: o_data_a = 16'b0000000000000000;
            14'h5e22: o_data_a = 16'b1111110010101000;
            14'h5e23: o_data_a = 16'b1111110000010000;
            14'h5e24: o_data_a = 16'b1110110010100000;
            14'h5e25: o_data_a = 16'b1111000010001000;
            14'h5e26: o_data_a = 16'b0000000000000000;
            14'h5e27: o_data_a = 16'b1111110010101000;
            14'h5e28: o_data_a = 16'b1111110000010000;
            14'h5e29: o_data_a = 16'b0000000000000001;
            14'h5e2a: o_data_a = 16'b1111110000100000;
            14'h5e2b: o_data_a = 16'b1110001100001000;
            14'h5e2c: o_data_a = 16'b0101110111011010;
            14'h5e2d: o_data_a = 16'b1110101010000111;
            14'h5e2e: o_data_a = 16'b0000000000000001;
            14'h5e2f: o_data_a = 16'b1111110000010000;
            14'h5e30: o_data_a = 16'b0000000000000011;
            14'h5e31: o_data_a = 16'b1110000010100000;
            14'h5e32: o_data_a = 16'b1111110000010000;
            14'h5e33: o_data_a = 16'b0000000000000000;
            14'h5e34: o_data_a = 16'b1111110111101000;
            14'h5e35: o_data_a = 16'b1110110010100000;
            14'h5e36: o_data_a = 16'b1110001100001000;
            14'h5e37: o_data_a = 16'b0000000000000001;
            14'h5e38: o_data_a = 16'b1111110000010000;
            14'h5e39: o_data_a = 16'b0000000000000100;
            14'h5e3a: o_data_a = 16'b1110000010100000;
            14'h5e3b: o_data_a = 16'b1111110000010000;
            14'h5e3c: o_data_a = 16'b0000000000000000;
            14'h5e3d: o_data_a = 16'b1111110111101000;
            14'h5e3e: o_data_a = 16'b1110110010100000;
            14'h5e3f: o_data_a = 16'b1110001100001000;
            14'h5e40: o_data_a = 16'b0000000000000010;
            14'h5e41: o_data_a = 16'b1110110000010000;
            14'h5e42: o_data_a = 16'b0000000000001101;
            14'h5e43: o_data_a = 16'b1110001100001000;
            14'h5e44: o_data_a = 16'b0101000011011101;
            14'h5e45: o_data_a = 16'b1110110000010000;
            14'h5e46: o_data_a = 16'b0000000000001110;
            14'h5e47: o_data_a = 16'b1110001100001000;
            14'h5e48: o_data_a = 16'b0101111001001100;
            14'h5e49: o_data_a = 16'b1110110000010000;
            14'h5e4a: o_data_a = 16'b0000000001011111;
            14'h5e4b: o_data_a = 16'b1110101010000111;
            14'h5e4c: o_data_a = 16'b0000000000000000;
            14'h5e4d: o_data_a = 16'b1111110010101000;
            14'h5e4e: o_data_a = 16'b1111110000010000;
            14'h5e4f: o_data_a = 16'b0000000000000101;
            14'h5e50: o_data_a = 16'b1110001100001000;
            14'h5e51: o_data_a = 16'b0000000000000000;
            14'h5e52: o_data_a = 16'b1111110111001000;
            14'h5e53: o_data_a = 16'b1111110010100000;
            14'h5e54: o_data_a = 16'b1110101010001000;
            14'h5e55: o_data_a = 16'b0000000000110110;
            14'h5e56: o_data_a = 16'b1110101010000111;
            14'h5e57: o_data_a = 16'b0000000000000010;
            14'h5e58: o_data_a = 16'b1111110111100000;
            14'h5e59: o_data_a = 16'b1111110000010000;
            14'h5e5a: o_data_a = 16'b0000000000000000;
            14'h5e5b: o_data_a = 16'b1111110111101000;
            14'h5e5c: o_data_a = 16'b1110110010100000;
            14'h5e5d: o_data_a = 16'b1110001100001000;
            14'h5e5e: o_data_a = 16'b0000000000000010;
            14'h5e5f: o_data_a = 16'b1111110000010000;
            14'h5e60: o_data_a = 16'b0000000000000011;
            14'h5e61: o_data_a = 16'b1110000010100000;
            14'h5e62: o_data_a = 16'b1111110000010000;
            14'h5e63: o_data_a = 16'b0000000000000000;
            14'h5e64: o_data_a = 16'b1111110111101000;
            14'h5e65: o_data_a = 16'b1110110010100000;
            14'h5e66: o_data_a = 16'b1110001100001000;
            14'h5e67: o_data_a = 16'b0000000000000000;
            14'h5e68: o_data_a = 16'b1111110010101000;
            14'h5e69: o_data_a = 16'b1111110000010000;
            14'h5e6a: o_data_a = 16'b1110110010100000;
            14'h5e6b: o_data_a = 16'b1111000111001000;
            14'h5e6c: o_data_a = 16'b0000000000000010;
            14'h5e6d: o_data_a = 16'b1111110000100000;
            14'h5e6e: o_data_a = 16'b1111110000010000;
            14'h5e6f: o_data_a = 16'b0000000000000000;
            14'h5e70: o_data_a = 16'b1111110111101000;
            14'h5e71: o_data_a = 16'b1110110010100000;
            14'h5e72: o_data_a = 16'b1110001100001000;
            14'h5e73: o_data_a = 16'b0000000000000010;
            14'h5e74: o_data_a = 16'b1111110111100000;
            14'h5e75: o_data_a = 16'b1110110111100000;
            14'h5e76: o_data_a = 16'b1111110000010000;
            14'h5e77: o_data_a = 16'b0000000000000000;
            14'h5e78: o_data_a = 16'b1111110111101000;
            14'h5e79: o_data_a = 16'b1110110010100000;
            14'h5e7a: o_data_a = 16'b1110001100001000;
            14'h5e7b: o_data_a = 16'b0000000000000000;
            14'h5e7c: o_data_a = 16'b1111110010101000;
            14'h5e7d: o_data_a = 16'b1111110000010000;
            14'h5e7e: o_data_a = 16'b1110110010100000;
            14'h5e7f: o_data_a = 16'b1111000010001000;
            14'h5e80: o_data_a = 16'b0000000000000010;
            14'h5e81: o_data_a = 16'b1111110000100000;
            14'h5e82: o_data_a = 16'b1111110000010000;
            14'h5e83: o_data_a = 16'b0000000000000000;
            14'h5e84: o_data_a = 16'b1111110111101000;
            14'h5e85: o_data_a = 16'b1110110010100000;
            14'h5e86: o_data_a = 16'b1110001100001000;
            14'h5e87: o_data_a = 16'b0000000000000010;
            14'h5e88: o_data_a = 16'b1111110111100000;
            14'h5e89: o_data_a = 16'b1110110111100000;
            14'h5e8a: o_data_a = 16'b1111110000010000;
            14'h5e8b: o_data_a = 16'b0000000000000000;
            14'h5e8c: o_data_a = 16'b1111110111101000;
            14'h5e8d: o_data_a = 16'b1110110010100000;
            14'h5e8e: o_data_a = 16'b1110001100001000;
            14'h5e8f: o_data_a = 16'b0000000000000000;
            14'h5e90: o_data_a = 16'b1111110010101000;
            14'h5e91: o_data_a = 16'b1111110000010000;
            14'h5e92: o_data_a = 16'b1110110010100000;
            14'h5e93: o_data_a = 16'b1111000111001000;
            14'h5e94: o_data_a = 16'b0000000000000011;
            14'h5e95: o_data_a = 16'b1110110000010000;
            14'h5e96: o_data_a = 16'b0000000000001101;
            14'h5e97: o_data_a = 16'b1110001100001000;
            14'h5e98: o_data_a = 16'b0101101011010011;
            14'h5e99: o_data_a = 16'b1110110000010000;
            14'h5e9a: o_data_a = 16'b0000000000001110;
            14'h5e9b: o_data_a = 16'b1110001100001000;
            14'h5e9c: o_data_a = 16'b0101111010100000;
            14'h5e9d: o_data_a = 16'b1110110000010000;
            14'h5e9e: o_data_a = 16'b0000000001011111;
            14'h5e9f: o_data_a = 16'b1110101010000111;
            14'h5ea0: o_data_a = 16'b0000000000000000;
            14'h5ea1: o_data_a = 16'b1111110010101000;
            14'h5ea2: o_data_a = 16'b1111110000010000;
            14'h5ea3: o_data_a = 16'b0000000000000101;
            14'h5ea4: o_data_a = 16'b1110001100001000;
            14'h5ea5: o_data_a = 16'b0000000000000010;
            14'h5ea6: o_data_a = 16'b1111110111100000;
            14'h5ea7: o_data_a = 16'b1111110000010000;
            14'h5ea8: o_data_a = 16'b0000000000000000;
            14'h5ea9: o_data_a = 16'b1111110111101000;
            14'h5eaa: o_data_a = 16'b1110110010100000;
            14'h5eab: o_data_a = 16'b1110001100001000;
            14'h5eac: o_data_a = 16'b0000000000000010;
            14'h5ead: o_data_a = 16'b1111110000010000;
            14'h5eae: o_data_a = 16'b0000000000000011;
            14'h5eaf: o_data_a = 16'b1110000010100000;
            14'h5eb0: o_data_a = 16'b1111110000010000;
            14'h5eb1: o_data_a = 16'b0000000000000000;
            14'h5eb2: o_data_a = 16'b1111110111101000;
            14'h5eb3: o_data_a = 16'b1110110010100000;
            14'h5eb4: o_data_a = 16'b1110001100001000;
            14'h5eb5: o_data_a = 16'b0000000000000000;
            14'h5eb6: o_data_a = 16'b1111110010101000;
            14'h5eb7: o_data_a = 16'b1111110000010000;
            14'h5eb8: o_data_a = 16'b1110110010100000;
            14'h5eb9: o_data_a = 16'b1111000010001000;
            14'h5eba: o_data_a = 16'b0000000000000010;
            14'h5ebb: o_data_a = 16'b1111110000100000;
            14'h5ebc: o_data_a = 16'b1111110000010000;
            14'h5ebd: o_data_a = 16'b0000000000000000;
            14'h5ebe: o_data_a = 16'b1111110111101000;
            14'h5ebf: o_data_a = 16'b1110110010100000;
            14'h5ec0: o_data_a = 16'b1110001100001000;
            14'h5ec1: o_data_a = 16'b0000000000000010;
            14'h5ec2: o_data_a = 16'b1111110111100000;
            14'h5ec3: o_data_a = 16'b1110110111100000;
            14'h5ec4: o_data_a = 16'b1111110000010000;
            14'h5ec5: o_data_a = 16'b0000000000000000;
            14'h5ec6: o_data_a = 16'b1111110111101000;
            14'h5ec7: o_data_a = 16'b1110110010100000;
            14'h5ec8: o_data_a = 16'b1110001100001000;
            14'h5ec9: o_data_a = 16'b0000000000000000;
            14'h5eca: o_data_a = 16'b1111110010101000;
            14'h5ecb: o_data_a = 16'b1111110000010000;
            14'h5ecc: o_data_a = 16'b1110110010100000;
            14'h5ecd: o_data_a = 16'b1111000010001000;
            14'h5ece: o_data_a = 16'b0000000000000010;
            14'h5ecf: o_data_a = 16'b1111110000100000;
            14'h5ed0: o_data_a = 16'b1111110000010000;
            14'h5ed1: o_data_a = 16'b0000000000000000;
            14'h5ed2: o_data_a = 16'b1111110111101000;
            14'h5ed3: o_data_a = 16'b1110110010100000;
            14'h5ed4: o_data_a = 16'b1110001100001000;
            14'h5ed5: o_data_a = 16'b0000000000000010;
            14'h5ed6: o_data_a = 16'b1111110111100000;
            14'h5ed7: o_data_a = 16'b1110110111100000;
            14'h5ed8: o_data_a = 16'b1111110000010000;
            14'h5ed9: o_data_a = 16'b0000000000000000;
            14'h5eda: o_data_a = 16'b1111110111101000;
            14'h5edb: o_data_a = 16'b1110110010100000;
            14'h5edc: o_data_a = 16'b1110001100001000;
            14'h5edd: o_data_a = 16'b0000000000000000;
            14'h5ede: o_data_a = 16'b1111110010101000;
            14'h5edf: o_data_a = 16'b1111110000010000;
            14'h5ee0: o_data_a = 16'b1110110010100000;
            14'h5ee1: o_data_a = 16'b1111000111001000;
            14'h5ee2: o_data_a = 16'b0000000000000011;
            14'h5ee3: o_data_a = 16'b1110110000010000;
            14'h5ee4: o_data_a = 16'b0000000000001101;
            14'h5ee5: o_data_a = 16'b1110001100001000;
            14'h5ee6: o_data_a = 16'b0101101011010011;
            14'h5ee7: o_data_a = 16'b1110110000010000;
            14'h5ee8: o_data_a = 16'b0000000000001110;
            14'h5ee9: o_data_a = 16'b1110001100001000;
            14'h5eea: o_data_a = 16'b0101111011101110;
            14'h5eeb: o_data_a = 16'b1110110000010000;
            14'h5eec: o_data_a = 16'b0000000001011111;
            14'h5eed: o_data_a = 16'b1110101010000111;
            14'h5eee: o_data_a = 16'b0000000000000000;
            14'h5eef: o_data_a = 16'b1111110010101000;
            14'h5ef0: o_data_a = 16'b1111110000010000;
            14'h5ef1: o_data_a = 16'b0000000000000101;
            14'h5ef2: o_data_a = 16'b1110001100001000;
            14'h5ef3: o_data_a = 16'b0000000000000010;
            14'h5ef4: o_data_a = 16'b1111110111100000;
            14'h5ef5: o_data_a = 16'b1111110000010000;
            14'h5ef6: o_data_a = 16'b0000000000000000;
            14'h5ef7: o_data_a = 16'b1111110111101000;
            14'h5ef8: o_data_a = 16'b1110110010100000;
            14'h5ef9: o_data_a = 16'b1110001100001000;
            14'h5efa: o_data_a = 16'b0000000000000010;
            14'h5efb: o_data_a = 16'b1111110111100000;
            14'h5efc: o_data_a = 16'b1110110111100000;
            14'h5efd: o_data_a = 16'b1111110000010000;
            14'h5efe: o_data_a = 16'b0000000000000000;
            14'h5eff: o_data_a = 16'b1111110111101000;
            14'h5f00: o_data_a = 16'b1110110010100000;
            14'h5f01: o_data_a = 16'b1110001100001000;
            14'h5f02: o_data_a = 16'b0000000000000000;
            14'h5f03: o_data_a = 16'b1111110010101000;
            14'h5f04: o_data_a = 16'b1111110000010000;
            14'h5f05: o_data_a = 16'b1110110010100000;
            14'h5f06: o_data_a = 16'b1111000111001000;
            14'h5f07: o_data_a = 16'b0000000000000010;
            14'h5f08: o_data_a = 16'b1111110000100000;
            14'h5f09: o_data_a = 16'b1111110000010000;
            14'h5f0a: o_data_a = 16'b0000000000000000;
            14'h5f0b: o_data_a = 16'b1111110111101000;
            14'h5f0c: o_data_a = 16'b1110110010100000;
            14'h5f0d: o_data_a = 16'b1110001100001000;
            14'h5f0e: o_data_a = 16'b0000000000000010;
            14'h5f0f: o_data_a = 16'b1111110000010000;
            14'h5f10: o_data_a = 16'b0000000000000011;
            14'h5f11: o_data_a = 16'b1110000010100000;
            14'h5f12: o_data_a = 16'b1111110000010000;
            14'h5f13: o_data_a = 16'b0000000000000000;
            14'h5f14: o_data_a = 16'b1111110111101000;
            14'h5f15: o_data_a = 16'b1110110010100000;
            14'h5f16: o_data_a = 16'b1110001100001000;
            14'h5f17: o_data_a = 16'b0000000000000000;
            14'h5f18: o_data_a = 16'b1111110010101000;
            14'h5f19: o_data_a = 16'b1111110000010000;
            14'h5f1a: o_data_a = 16'b1110110010100000;
            14'h5f1b: o_data_a = 16'b1111000111001000;
            14'h5f1c: o_data_a = 16'b0000000000000010;
            14'h5f1d: o_data_a = 16'b1111110000100000;
            14'h5f1e: o_data_a = 16'b1111110000010000;
            14'h5f1f: o_data_a = 16'b0000000000000000;
            14'h5f20: o_data_a = 16'b1111110111101000;
            14'h5f21: o_data_a = 16'b1110110010100000;
            14'h5f22: o_data_a = 16'b1110001100001000;
            14'h5f23: o_data_a = 16'b0000000000000010;
            14'h5f24: o_data_a = 16'b1111110000010000;
            14'h5f25: o_data_a = 16'b0000000000000011;
            14'h5f26: o_data_a = 16'b1110000010100000;
            14'h5f27: o_data_a = 16'b1111110000010000;
            14'h5f28: o_data_a = 16'b0000000000000000;
            14'h5f29: o_data_a = 16'b1111110111101000;
            14'h5f2a: o_data_a = 16'b1110110010100000;
            14'h5f2b: o_data_a = 16'b1110001100001000;
            14'h5f2c: o_data_a = 16'b0000000000000000;
            14'h5f2d: o_data_a = 16'b1111110010101000;
            14'h5f2e: o_data_a = 16'b1111110000010000;
            14'h5f2f: o_data_a = 16'b1110110010100000;
            14'h5f30: o_data_a = 16'b1111000010001000;
            14'h5f31: o_data_a = 16'b0000000000000011;
            14'h5f32: o_data_a = 16'b1110110000010000;
            14'h5f33: o_data_a = 16'b0000000000001101;
            14'h5f34: o_data_a = 16'b1110001100001000;
            14'h5f35: o_data_a = 16'b0101101011010011;
            14'h5f36: o_data_a = 16'b1110110000010000;
            14'h5f37: o_data_a = 16'b0000000000001110;
            14'h5f38: o_data_a = 16'b1110001100001000;
            14'h5f39: o_data_a = 16'b0101111100111101;
            14'h5f3a: o_data_a = 16'b1110110000010000;
            14'h5f3b: o_data_a = 16'b0000000001011111;
            14'h5f3c: o_data_a = 16'b1110101010000111;
            14'h5f3d: o_data_a = 16'b0000000000000000;
            14'h5f3e: o_data_a = 16'b1111110010101000;
            14'h5f3f: o_data_a = 16'b1111110000010000;
            14'h5f40: o_data_a = 16'b0000000000000101;
            14'h5f41: o_data_a = 16'b1110001100001000;
            14'h5f42: o_data_a = 16'b0000000000000010;
            14'h5f43: o_data_a = 16'b1111110111100000;
            14'h5f44: o_data_a = 16'b1111110000010000;
            14'h5f45: o_data_a = 16'b0000000000000000;
            14'h5f46: o_data_a = 16'b1111110111101000;
            14'h5f47: o_data_a = 16'b1110110010100000;
            14'h5f48: o_data_a = 16'b1110001100001000;
            14'h5f49: o_data_a = 16'b0000000000000010;
            14'h5f4a: o_data_a = 16'b1111110111100000;
            14'h5f4b: o_data_a = 16'b1110110111100000;
            14'h5f4c: o_data_a = 16'b1111110000010000;
            14'h5f4d: o_data_a = 16'b0000000000000000;
            14'h5f4e: o_data_a = 16'b1111110111101000;
            14'h5f4f: o_data_a = 16'b1110110010100000;
            14'h5f50: o_data_a = 16'b1110001100001000;
            14'h5f51: o_data_a = 16'b0000000000000000;
            14'h5f52: o_data_a = 16'b1111110010101000;
            14'h5f53: o_data_a = 16'b1111110000010000;
            14'h5f54: o_data_a = 16'b1110110010100000;
            14'h5f55: o_data_a = 16'b1111000010001000;
            14'h5f56: o_data_a = 16'b0000000000000010;
            14'h5f57: o_data_a = 16'b1111110000100000;
            14'h5f58: o_data_a = 16'b1111110000010000;
            14'h5f59: o_data_a = 16'b0000000000000000;
            14'h5f5a: o_data_a = 16'b1111110111101000;
            14'h5f5b: o_data_a = 16'b1110110010100000;
            14'h5f5c: o_data_a = 16'b1110001100001000;
            14'h5f5d: o_data_a = 16'b0000000000000010;
            14'h5f5e: o_data_a = 16'b1111110000010000;
            14'h5f5f: o_data_a = 16'b0000000000000011;
            14'h5f60: o_data_a = 16'b1110000010100000;
            14'h5f61: o_data_a = 16'b1111110000010000;
            14'h5f62: o_data_a = 16'b0000000000000000;
            14'h5f63: o_data_a = 16'b1111110111101000;
            14'h5f64: o_data_a = 16'b1110110010100000;
            14'h5f65: o_data_a = 16'b1110001100001000;
            14'h5f66: o_data_a = 16'b0000000000000000;
            14'h5f67: o_data_a = 16'b1111110010101000;
            14'h5f68: o_data_a = 16'b1111110000010000;
            14'h5f69: o_data_a = 16'b1110110010100000;
            14'h5f6a: o_data_a = 16'b1111000111001000;
            14'h5f6b: o_data_a = 16'b0000000000000010;
            14'h5f6c: o_data_a = 16'b1111110000100000;
            14'h5f6d: o_data_a = 16'b1111110000010000;
            14'h5f6e: o_data_a = 16'b0000000000000000;
            14'h5f6f: o_data_a = 16'b1111110111101000;
            14'h5f70: o_data_a = 16'b1110110010100000;
            14'h5f71: o_data_a = 16'b1110001100001000;
            14'h5f72: o_data_a = 16'b0000000000000010;
            14'h5f73: o_data_a = 16'b1111110000010000;
            14'h5f74: o_data_a = 16'b0000000000000011;
            14'h5f75: o_data_a = 16'b1110000010100000;
            14'h5f76: o_data_a = 16'b1111110000010000;
            14'h5f77: o_data_a = 16'b0000000000000000;
            14'h5f78: o_data_a = 16'b1111110111101000;
            14'h5f79: o_data_a = 16'b1110110010100000;
            14'h5f7a: o_data_a = 16'b1110001100001000;
            14'h5f7b: o_data_a = 16'b0000000000000000;
            14'h5f7c: o_data_a = 16'b1111110010101000;
            14'h5f7d: o_data_a = 16'b1111110000010000;
            14'h5f7e: o_data_a = 16'b1110110010100000;
            14'h5f7f: o_data_a = 16'b1111000010001000;
            14'h5f80: o_data_a = 16'b0000000000000011;
            14'h5f81: o_data_a = 16'b1110110000010000;
            14'h5f82: o_data_a = 16'b0000000000001101;
            14'h5f83: o_data_a = 16'b1110001100001000;
            14'h5f84: o_data_a = 16'b0101101011010011;
            14'h5f85: o_data_a = 16'b1110110000010000;
            14'h5f86: o_data_a = 16'b0000000000001110;
            14'h5f87: o_data_a = 16'b1110001100001000;
            14'h5f88: o_data_a = 16'b0101111110001100;
            14'h5f89: o_data_a = 16'b1110110000010000;
            14'h5f8a: o_data_a = 16'b0000000001011111;
            14'h5f8b: o_data_a = 16'b1110101010000111;
            14'h5f8c: o_data_a = 16'b0000000000000000;
            14'h5f8d: o_data_a = 16'b1111110010101000;
            14'h5f8e: o_data_a = 16'b1111110000010000;
            14'h5f8f: o_data_a = 16'b0000000000000101;
            14'h5f90: o_data_a = 16'b1110001100001000;
            14'h5f91: o_data_a = 16'b0000000000000000;
            14'h5f92: o_data_a = 16'b1111110111001000;
            14'h5f93: o_data_a = 16'b1111110010100000;
            14'h5f94: o_data_a = 16'b1110101010001000;
            14'h5f95: o_data_a = 16'b0000000000110110;
            14'h5f96: o_data_a = 16'b1110101010000111;
            14'h5f97: o_data_a = 16'b0000000000000011;
            14'h5f98: o_data_a = 16'b1110110000010000;
            14'h5f99: o_data_a = 16'b1110001110010000;
            14'h5f9a: o_data_a = 16'b0000000000000000;
            14'h5f9b: o_data_a = 16'b1111110111101000;
            14'h5f9c: o_data_a = 16'b1110110010100000;
            14'h5f9d: o_data_a = 16'b1110101010001000;
            14'h5f9e: o_data_a = 16'b0101111110011001;
            14'h5f9f: o_data_a = 16'b1110001100000001;
            14'h5fa0: o_data_a = 16'b0000000000000010;
            14'h5fa1: o_data_a = 16'b1111110000100000;
            14'h5fa2: o_data_a = 16'b1111110000010000;
            14'h5fa3: o_data_a = 16'b0000000000000000;
            14'h5fa4: o_data_a = 16'b1111110111101000;
            14'h5fa5: o_data_a = 16'b1110110010100000;
            14'h5fa6: o_data_a = 16'b1110001100001000;
            14'h5fa7: o_data_a = 16'b0000000000000000;
            14'h5fa8: o_data_a = 16'b1111110111001000;
            14'h5fa9: o_data_a = 16'b1111110010100000;
            14'h5faa: o_data_a = 16'b1110101010001000;
            14'h5fab: o_data_a = 16'b0101111110101111;
            14'h5fac: o_data_a = 16'b1110110000010000;
            14'h5fad: o_data_a = 16'b0000000000100110;
            14'h5fae: o_data_a = 16'b1110101010000111;
            14'h5faf: o_data_a = 16'b0000000000000010;
            14'h5fb0: o_data_a = 16'b1111110000100000;
            14'h5fb1: o_data_a = 16'b1111110000010000;
            14'h5fb2: o_data_a = 16'b0000000000000000;
            14'h5fb3: o_data_a = 16'b1111110111101000;
            14'h5fb4: o_data_a = 16'b1110110010100000;
            14'h5fb5: o_data_a = 16'b1110001100001000;
            14'h5fb6: o_data_a = 16'b0000000111111111;
            14'h5fb7: o_data_a = 16'b1110110000010000;
            14'h5fb8: o_data_a = 16'b0000000000000000;
            14'h5fb9: o_data_a = 16'b1111110111101000;
            14'h5fba: o_data_a = 16'b1110110010100000;
            14'h5fbb: o_data_a = 16'b1110001100001000;
            14'h5fbc: o_data_a = 16'b0101111111000000;
            14'h5fbd: o_data_a = 16'b1110110000010000;
            14'h5fbe: o_data_a = 16'b0000000000010110;
            14'h5fbf: o_data_a = 16'b1110101010000111;
            14'h5fc0: o_data_a = 16'b0000000000000000;
            14'h5fc1: o_data_a = 16'b1111110010101000;
            14'h5fc2: o_data_a = 16'b1111110000010000;
            14'h5fc3: o_data_a = 16'b1110110010100000;
            14'h5fc4: o_data_a = 16'b1111010101001000;
            14'h5fc5: o_data_a = 16'b0000000000000010;
            14'h5fc6: o_data_a = 16'b1111110111100000;
            14'h5fc7: o_data_a = 16'b1111110000010000;
            14'h5fc8: o_data_a = 16'b0000000000000000;
            14'h5fc9: o_data_a = 16'b1111110111101000;
            14'h5fca: o_data_a = 16'b1110110010100000;
            14'h5fcb: o_data_a = 16'b1110001100001000;
            14'h5fcc: o_data_a = 16'b0000000000000000;
            14'h5fcd: o_data_a = 16'b1111110111001000;
            14'h5fce: o_data_a = 16'b1111110010100000;
            14'h5fcf: o_data_a = 16'b1110101010001000;
            14'h5fd0: o_data_a = 16'b0101111111010100;
            14'h5fd1: o_data_a = 16'b1110110000010000;
            14'h5fd2: o_data_a = 16'b0000000000100110;
            14'h5fd3: o_data_a = 16'b1110101010000111;
            14'h5fd4: o_data_a = 16'b0000000000000000;
            14'h5fd5: o_data_a = 16'b1111110010101000;
            14'h5fd6: o_data_a = 16'b1111110000010000;
            14'h5fd7: o_data_a = 16'b1110110010100000;
            14'h5fd8: o_data_a = 16'b1111010101001000;
            14'h5fd9: o_data_a = 16'b0000000000000010;
            14'h5fda: o_data_a = 16'b1111110111100000;
            14'h5fdb: o_data_a = 16'b1111110000010000;
            14'h5fdc: o_data_a = 16'b0000000000000000;
            14'h5fdd: o_data_a = 16'b1111110111101000;
            14'h5fde: o_data_a = 16'b1110110010100000;
            14'h5fdf: o_data_a = 16'b1110001100001000;
            14'h5fe0: o_data_a = 16'b0000000011111111;
            14'h5fe1: o_data_a = 16'b1110110000010000;
            14'h5fe2: o_data_a = 16'b0000000000000000;
            14'h5fe3: o_data_a = 16'b1111110111101000;
            14'h5fe4: o_data_a = 16'b1110110010100000;
            14'h5fe5: o_data_a = 16'b1110001100001000;
            14'h5fe6: o_data_a = 16'b0101111111101010;
            14'h5fe7: o_data_a = 16'b1110110000010000;
            14'h5fe8: o_data_a = 16'b0000000000010110;
            14'h5fe9: o_data_a = 16'b1110101010000111;
            14'h5fea: o_data_a = 16'b0000000000000000;
            14'h5feb: o_data_a = 16'b1111110010101000;
            14'h5fec: o_data_a = 16'b1111110000010000;
            14'h5fed: o_data_a = 16'b1110110010100000;
            14'h5fee: o_data_a = 16'b1111010101001000;
            14'h5fef: o_data_a = 16'b0000000000000000;
            14'h5ff0: o_data_a = 16'b1111110010101000;
            14'h5ff1: o_data_a = 16'b1111110000010000;
            14'h5ff2: o_data_a = 16'b0101111111110110;
            14'h5ff3: o_data_a = 16'b1110001100000101;
            14'h5ff4: o_data_a = 16'b0110000000001101;
            14'h5ff5: o_data_a = 16'b1110101010000111;
            14'h5ff6: o_data_a = 16'b0000000000001100;
            14'h5ff7: o_data_a = 16'b1110110000010000;
            14'h5ff8: o_data_a = 16'b0000000000000000;
            14'h5ff9: o_data_a = 16'b1111110111101000;
            14'h5ffa: o_data_a = 16'b1110110010100000;
            14'h5ffb: o_data_a = 16'b1110001100001000;
            14'h5ffc: o_data_a = 16'b0000000000000001;
            14'h5ffd: o_data_a = 16'b1110110000010000;
            14'h5ffe: o_data_a = 16'b0000000000001101;
            14'h5fff: o_data_a = 16'b1110001100001000;
            14'h6000: o_data_a = 16'b0110101011011001;
            14'h6001: o_data_a = 16'b1110110000010000;
            14'h6002: o_data_a = 16'b0000000000001110;
            14'h6003: o_data_a = 16'b1110001100001000;
            14'h6004: o_data_a = 16'b0110000000001000;
            14'h6005: o_data_a = 16'b1110110000010000;
            14'h6006: o_data_a = 16'b0000000001011111;
            14'h6007: o_data_a = 16'b1110101010000111;
            14'h6008: o_data_a = 16'b0000000000000000;
            14'h6009: o_data_a = 16'b1111110010101000;
            14'h600a: o_data_a = 16'b1111110000010000;
            14'h600b: o_data_a = 16'b0000000000000101;
            14'h600c: o_data_a = 16'b1110001100001000;
            14'h600d: o_data_a = 16'b0000000000000010;
            14'h600e: o_data_a = 16'b1111110000100000;
            14'h600f: o_data_a = 16'b1111110000010000;
            14'h6010: o_data_a = 16'b0000000000000000;
            14'h6011: o_data_a = 16'b1111110111101000;
            14'h6012: o_data_a = 16'b1110110010100000;
            14'h6013: o_data_a = 16'b1110001100001000;
            14'h6014: o_data_a = 16'b0000000000000010;
            14'h6015: o_data_a = 16'b1111110111100000;
            14'h6016: o_data_a = 16'b1110110111100000;
            14'h6017: o_data_a = 16'b1111110000010000;
            14'h6018: o_data_a = 16'b0000000000000000;
            14'h6019: o_data_a = 16'b1111110111101000;
            14'h601a: o_data_a = 16'b1110110010100000;
            14'h601b: o_data_a = 16'b1110001100001000;
            14'h601c: o_data_a = 16'b0000000000000000;
            14'h601d: o_data_a = 16'b1111110010101000;
            14'h601e: o_data_a = 16'b1111110000010000;
            14'h601f: o_data_a = 16'b1110110010100000;
            14'h6020: o_data_a = 16'b1111000111001000;
            14'h6021: o_data_a = 16'b0000000000000000;
            14'h6022: o_data_a = 16'b1111110111001000;
            14'h6023: o_data_a = 16'b1111110010100000;
            14'h6024: o_data_a = 16'b1110101010001000;
            14'h6025: o_data_a = 16'b0110000000101001;
            14'h6026: o_data_a = 16'b1110110000010000;
            14'h6027: o_data_a = 16'b0000000000100110;
            14'h6028: o_data_a = 16'b1110101010000111;
            14'h6029: o_data_a = 16'b0000000000000010;
            14'h602a: o_data_a = 16'b1111110000100000;
            14'h602b: o_data_a = 16'b1111110000010000;
            14'h602c: o_data_a = 16'b0000000000000000;
            14'h602d: o_data_a = 16'b1111110111101000;
            14'h602e: o_data_a = 16'b1110110010100000;
            14'h602f: o_data_a = 16'b1110001100001000;
            14'h6030: o_data_a = 16'b0000000000000010;
            14'h6031: o_data_a = 16'b1111110111100000;
            14'h6032: o_data_a = 16'b1110110111100000;
            14'h6033: o_data_a = 16'b1111110000010000;
            14'h6034: o_data_a = 16'b0000000000000000;
            14'h6035: o_data_a = 16'b1111110111101000;
            14'h6036: o_data_a = 16'b1110110010100000;
            14'h6037: o_data_a = 16'b1110001100001000;
            14'h6038: o_data_a = 16'b0000000000000000;
            14'h6039: o_data_a = 16'b1111110010101000;
            14'h603a: o_data_a = 16'b1111110000010000;
            14'h603b: o_data_a = 16'b1110110010100000;
            14'h603c: o_data_a = 16'b1111000010001000;
            14'h603d: o_data_a = 16'b0000000111111111;
            14'h603e: o_data_a = 16'b1110110000010000;
            14'h603f: o_data_a = 16'b0000000000000000;
            14'h6040: o_data_a = 16'b1111110111101000;
            14'h6041: o_data_a = 16'b1110110010100000;
            14'h6042: o_data_a = 16'b1110001100001000;
            14'h6043: o_data_a = 16'b0110000001000111;
            14'h6044: o_data_a = 16'b1110110000010000;
            14'h6045: o_data_a = 16'b0000000000010110;
            14'h6046: o_data_a = 16'b1110101010000111;
            14'h6047: o_data_a = 16'b0000000000000000;
            14'h6048: o_data_a = 16'b1111110010101000;
            14'h6049: o_data_a = 16'b1111110000010000;
            14'h604a: o_data_a = 16'b1110110010100000;
            14'h604b: o_data_a = 16'b1111010101001000;
            14'h604c: o_data_a = 16'b0000000000000010;
            14'h604d: o_data_a = 16'b1111110111100000;
            14'h604e: o_data_a = 16'b1111110000010000;
            14'h604f: o_data_a = 16'b0000000000000000;
            14'h6050: o_data_a = 16'b1111110111101000;
            14'h6051: o_data_a = 16'b1110110010100000;
            14'h6052: o_data_a = 16'b1110001100001000;
            14'h6053: o_data_a = 16'b0000000000000010;
            14'h6054: o_data_a = 16'b1111110111100000;
            14'h6055: o_data_a = 16'b1110110111100000;
            14'h6056: o_data_a = 16'b1111110000010000;
            14'h6057: o_data_a = 16'b0000000000000000;
            14'h6058: o_data_a = 16'b1111110111101000;
            14'h6059: o_data_a = 16'b1110110010100000;
            14'h605a: o_data_a = 16'b1110001100001000;
            14'h605b: o_data_a = 16'b0000000000000000;
            14'h605c: o_data_a = 16'b1111110010101000;
            14'h605d: o_data_a = 16'b1111110000010000;
            14'h605e: o_data_a = 16'b1110110010100000;
            14'h605f: o_data_a = 16'b1111000111001000;
            14'h6060: o_data_a = 16'b0000000000000000;
            14'h6061: o_data_a = 16'b1111110111001000;
            14'h6062: o_data_a = 16'b1111110010100000;
            14'h6063: o_data_a = 16'b1110101010001000;
            14'h6064: o_data_a = 16'b0110000001101000;
            14'h6065: o_data_a = 16'b1110110000010000;
            14'h6066: o_data_a = 16'b0000000000100110;
            14'h6067: o_data_a = 16'b1110101010000111;
            14'h6068: o_data_a = 16'b0000000000000000;
            14'h6069: o_data_a = 16'b1111110010101000;
            14'h606a: o_data_a = 16'b1111110000010000;
            14'h606b: o_data_a = 16'b1110110010100000;
            14'h606c: o_data_a = 16'b1111010101001000;
            14'h606d: o_data_a = 16'b0000000000000010;
            14'h606e: o_data_a = 16'b1111110111100000;
            14'h606f: o_data_a = 16'b1111110000010000;
            14'h6070: o_data_a = 16'b0000000000000000;
            14'h6071: o_data_a = 16'b1111110111101000;
            14'h6072: o_data_a = 16'b1110110010100000;
            14'h6073: o_data_a = 16'b1110001100001000;
            14'h6074: o_data_a = 16'b0000000000000010;
            14'h6075: o_data_a = 16'b1111110111100000;
            14'h6076: o_data_a = 16'b1110110111100000;
            14'h6077: o_data_a = 16'b1111110000010000;
            14'h6078: o_data_a = 16'b0000000000000000;
            14'h6079: o_data_a = 16'b1111110111101000;
            14'h607a: o_data_a = 16'b1110110010100000;
            14'h607b: o_data_a = 16'b1110001100001000;
            14'h607c: o_data_a = 16'b0000000000000000;
            14'h607d: o_data_a = 16'b1111110010101000;
            14'h607e: o_data_a = 16'b1111110000010000;
            14'h607f: o_data_a = 16'b1110110010100000;
            14'h6080: o_data_a = 16'b1111000010001000;
            14'h6081: o_data_a = 16'b0000000011111111;
            14'h6082: o_data_a = 16'b1110110000010000;
            14'h6083: o_data_a = 16'b0000000000000000;
            14'h6084: o_data_a = 16'b1111110111101000;
            14'h6085: o_data_a = 16'b1110110010100000;
            14'h6086: o_data_a = 16'b1110001100001000;
            14'h6087: o_data_a = 16'b0110000010001011;
            14'h6088: o_data_a = 16'b1110110000010000;
            14'h6089: o_data_a = 16'b0000000000010110;
            14'h608a: o_data_a = 16'b1110101010000111;
            14'h608b: o_data_a = 16'b0000000000000000;
            14'h608c: o_data_a = 16'b1111110010101000;
            14'h608d: o_data_a = 16'b1111110000010000;
            14'h608e: o_data_a = 16'b1110110010100000;
            14'h608f: o_data_a = 16'b1111010101001000;
            14'h6090: o_data_a = 16'b0000000000000000;
            14'h6091: o_data_a = 16'b1111110010101000;
            14'h6092: o_data_a = 16'b1111110000010000;
            14'h6093: o_data_a = 16'b0110000010010111;
            14'h6094: o_data_a = 16'b1110001100000101;
            14'h6095: o_data_a = 16'b0110000010101110;
            14'h6096: o_data_a = 16'b1110101010000111;
            14'h6097: o_data_a = 16'b0000000000001101;
            14'h6098: o_data_a = 16'b1110110000010000;
            14'h6099: o_data_a = 16'b0000000000000000;
            14'h609a: o_data_a = 16'b1111110111101000;
            14'h609b: o_data_a = 16'b1110110010100000;
            14'h609c: o_data_a = 16'b1110001100001000;
            14'h609d: o_data_a = 16'b0000000000000001;
            14'h609e: o_data_a = 16'b1110110000010000;
            14'h609f: o_data_a = 16'b0000000000001101;
            14'h60a0: o_data_a = 16'b1110001100001000;
            14'h60a1: o_data_a = 16'b0110101011011001;
            14'h60a2: o_data_a = 16'b1110110000010000;
            14'h60a3: o_data_a = 16'b0000000000001110;
            14'h60a4: o_data_a = 16'b1110001100001000;
            14'h60a5: o_data_a = 16'b0110000010101001;
            14'h60a6: o_data_a = 16'b1110110000010000;
            14'h60a7: o_data_a = 16'b0000000001011111;
            14'h60a8: o_data_a = 16'b1110101010000111;
            14'h60a9: o_data_a = 16'b0000000000000000;
            14'h60aa: o_data_a = 16'b1111110010101000;
            14'h60ab: o_data_a = 16'b1111110000010000;
            14'h60ac: o_data_a = 16'b0000000000000101;
            14'h60ad: o_data_a = 16'b1110001100001000;
            14'h60ae: o_data_a = 16'b0000000000000010;
            14'h60af: o_data_a = 16'b1111110111100000;
            14'h60b0: o_data_a = 16'b1110110111100000;
            14'h60b1: o_data_a = 16'b1111110000010000;
            14'h60b2: o_data_a = 16'b0000000000000000;
            14'h60b3: o_data_a = 16'b1111110111101000;
            14'h60b4: o_data_a = 16'b1110110010100000;
            14'h60b5: o_data_a = 16'b1110001100001000;
            14'h60b6: o_data_a = 16'b0000000000000000;
            14'h60b7: o_data_a = 16'b1111110010101000;
            14'h60b8: o_data_a = 16'b1111110000010000;
            14'h60b9: o_data_a = 16'b0000000000000001;
            14'h60ba: o_data_a = 16'b1111110111100000;
            14'h60bb: o_data_a = 16'b1110001100001000;
            14'h60bc: o_data_a = 16'b0000000000000000;
            14'h60bd: o_data_a = 16'b1111110111001000;
            14'h60be: o_data_a = 16'b1111110010100000;
            14'h60bf: o_data_a = 16'b1110111111001000;
            14'h60c0: o_data_a = 16'b0000000000000010;
            14'h60c1: o_data_a = 16'b1111110111100000;
            14'h60c2: o_data_a = 16'b1110110111100000;
            14'h60c3: o_data_a = 16'b1111110000010000;
            14'h60c4: o_data_a = 16'b0000000000000000;
            14'h60c5: o_data_a = 16'b1111110111101000;
            14'h60c6: o_data_a = 16'b1110110010100000;
            14'h60c7: o_data_a = 16'b1110001100001000;
            14'h60c8: o_data_a = 16'b0000000000000000;
            14'h60c9: o_data_a = 16'b1111110010101000;
            14'h60ca: o_data_a = 16'b1111110000010000;
            14'h60cb: o_data_a = 16'b1110110010100000;
            14'h60cc: o_data_a = 16'b1111000111001000;
            14'h60cd: o_data_a = 16'b0000000000000000;
            14'h60ce: o_data_a = 16'b1111110010101000;
            14'h60cf: o_data_a = 16'b1111110000010000;
            14'h60d0: o_data_a = 16'b0000000000000001;
            14'h60d1: o_data_a = 16'b1111110111100000;
            14'h60d2: o_data_a = 16'b1110110111100000;
            14'h60d3: o_data_a = 16'b1110001100001000;
            14'h60d4: o_data_a = 16'b0000000000000010;
            14'h60d5: o_data_a = 16'b1111110000100000;
            14'h60d6: o_data_a = 16'b1111110000010000;
            14'h60d7: o_data_a = 16'b0000000000000000;
            14'h60d8: o_data_a = 16'b1111110111101000;
            14'h60d9: o_data_a = 16'b1110110010100000;
            14'h60da: o_data_a = 16'b1110001100001000;
            14'h60db: o_data_a = 16'b0000000000000010;
            14'h60dc: o_data_a = 16'b1111110111100000;
            14'h60dd: o_data_a = 16'b1111110000010000;
            14'h60de: o_data_a = 16'b0000000000000000;
            14'h60df: o_data_a = 16'b1111110111101000;
            14'h60e0: o_data_a = 16'b1110110010100000;
            14'h60e1: o_data_a = 16'b1110001100001000;
            14'h60e2: o_data_a = 16'b0000000000000001;
            14'h60e3: o_data_a = 16'b1111110000100000;
            14'h60e4: o_data_a = 16'b1111110000010000;
            14'h60e5: o_data_a = 16'b0000000000000000;
            14'h60e6: o_data_a = 16'b1111110111101000;
            14'h60e7: o_data_a = 16'b1110110010100000;
            14'h60e8: o_data_a = 16'b1110001100001000;
            14'h60e9: o_data_a = 16'b0000000000000001;
            14'h60ea: o_data_a = 16'b1111110111100000;
            14'h60eb: o_data_a = 16'b1111110000010000;
            14'h60ec: o_data_a = 16'b0000000000000000;
            14'h60ed: o_data_a = 16'b1111110111101000;
            14'h60ee: o_data_a = 16'b1110110010100000;
            14'h60ef: o_data_a = 16'b1110001100001000;
            14'h60f0: o_data_a = 16'b0000000000000100;
            14'h60f1: o_data_a = 16'b1110110000010000;
            14'h60f2: o_data_a = 16'b0000000000001101;
            14'h60f3: o_data_a = 16'b1110001100001000;
            14'h60f4: o_data_a = 16'b0101111001010111;
            14'h60f5: o_data_a = 16'b1110110000010000;
            14'h60f6: o_data_a = 16'b0000000000001110;
            14'h60f7: o_data_a = 16'b1110001100001000;
            14'h60f8: o_data_a = 16'b0110000011111100;
            14'h60f9: o_data_a = 16'b1110110000010000;
            14'h60fa: o_data_a = 16'b0000000001011111;
            14'h60fb: o_data_a = 16'b1110101010000111;
            14'h60fc: o_data_a = 16'b0000000000000000;
            14'h60fd: o_data_a = 16'b1111110010101000;
            14'h60fe: o_data_a = 16'b1111110000010000;
            14'h60ff: o_data_a = 16'b0000000000000101;
            14'h6100: o_data_a = 16'b1110001100001000;
            14'h6101: o_data_a = 16'b0000000000000001;
            14'h6102: o_data_a = 16'b1111110111100000;
            14'h6103: o_data_a = 16'b1111110000010000;
            14'h6104: o_data_a = 16'b0000000000000000;
            14'h6105: o_data_a = 16'b1111110111101000;
            14'h6106: o_data_a = 16'b1110110010100000;
            14'h6107: o_data_a = 16'b1110001100001000;
            14'h6108: o_data_a = 16'b0000000000000001;
            14'h6109: o_data_a = 16'b1111110000100000;
            14'h610a: o_data_a = 16'b1111110000010000;
            14'h610b: o_data_a = 16'b0000000000000000;
            14'h610c: o_data_a = 16'b1111110111101000;
            14'h610d: o_data_a = 16'b1110110010100000;
            14'h610e: o_data_a = 16'b1110001100001000;
            14'h610f: o_data_a = 16'b0110000100010011;
            14'h6110: o_data_a = 16'b1110110000010000;
            14'h6111: o_data_a = 16'b0000000000010110;
            14'h6112: o_data_a = 16'b1110101010000111;
            14'h6113: o_data_a = 16'b0000000000000000;
            14'h6114: o_data_a = 16'b1111110010100000;
            14'h6115: o_data_a = 16'b1111110001001000;
            14'h6116: o_data_a = 16'b0000000000000000;
            14'h6117: o_data_a = 16'b1111110010101000;
            14'h6118: o_data_a = 16'b1111110000010000;
            14'h6119: o_data_a = 16'b0110001000001011;
            14'h611a: o_data_a = 16'b1110001100000101;
            14'h611b: o_data_a = 16'b0000000000000001;
            14'h611c: o_data_a = 16'b1111110111100000;
            14'h611d: o_data_a = 16'b1110110111100000;
            14'h611e: o_data_a = 16'b1111110000010000;
            14'h611f: o_data_a = 16'b0000000000000000;
            14'h6120: o_data_a = 16'b1111110111101000;
            14'h6121: o_data_a = 16'b1110110010100000;
            14'h6122: o_data_a = 16'b1110001100001000;
            14'h6123: o_data_a = 16'b0000000000000000;
            14'h6124: o_data_a = 16'b1111110111001000;
            14'h6125: o_data_a = 16'b1111110010100000;
            14'h6126: o_data_a = 16'b1110101010001000;
            14'h6127: o_data_a = 16'b0110000100101011;
            14'h6128: o_data_a = 16'b1110110000010000;
            14'h6129: o_data_a = 16'b0000000000100110;
            14'h612a: o_data_a = 16'b1110101010000111;
            14'h612b: o_data_a = 16'b0000000000000000;
            14'h612c: o_data_a = 16'b1111110010101000;
            14'h612d: o_data_a = 16'b1111110000010000;
            14'h612e: o_data_a = 16'b0110000100110010;
            14'h612f: o_data_a = 16'b1110001100000101;
            14'h6130: o_data_a = 16'b0110000101101100;
            14'h6131: o_data_a = 16'b1110101010000111;
            14'h6132: o_data_a = 16'b0000000000000001;
            14'h6133: o_data_a = 16'b1111110111100000;
            14'h6134: o_data_a = 16'b1110110111100000;
            14'h6135: o_data_a = 16'b1111110000010000;
            14'h6136: o_data_a = 16'b0000000000000000;
            14'h6137: o_data_a = 16'b1111110111101000;
            14'h6138: o_data_a = 16'b1110110010100000;
            14'h6139: o_data_a = 16'b1110001100001000;
            14'h613a: o_data_a = 16'b0000000000000010;
            14'h613b: o_data_a = 16'b1110110000010000;
            14'h613c: o_data_a = 16'b0000000000000000;
            14'h613d: o_data_a = 16'b1111110111101000;
            14'h613e: o_data_a = 16'b1110110010100000;
            14'h613f: o_data_a = 16'b1110001100001000;
            14'h6140: o_data_a = 16'b0000000000000001;
            14'h6141: o_data_a = 16'b1111110000100000;
            14'h6142: o_data_a = 16'b1111110000010000;
            14'h6143: o_data_a = 16'b0000000000000000;
            14'h6144: o_data_a = 16'b1111110111101000;
            14'h6145: o_data_a = 16'b1110110010100000;
            14'h6146: o_data_a = 16'b1110001100001000;
            14'h6147: o_data_a = 16'b0000000000000010;
            14'h6148: o_data_a = 16'b1110110000010000;
            14'h6149: o_data_a = 16'b0000000000001101;
            14'h614a: o_data_a = 16'b1110001100001000;
            14'h614b: o_data_a = 16'b0001101010100110;
            14'h614c: o_data_a = 16'b1110110000010000;
            14'h614d: o_data_a = 16'b0000000000001110;
            14'h614e: o_data_a = 16'b1110001100001000;
            14'h614f: o_data_a = 16'b0110000101010011;
            14'h6150: o_data_a = 16'b1110110000010000;
            14'h6151: o_data_a = 16'b0000000001011111;
            14'h6152: o_data_a = 16'b1110101010000111;
            14'h6153: o_data_a = 16'b0000000000000000;
            14'h6154: o_data_a = 16'b1111110010101000;
            14'h6155: o_data_a = 16'b1111110000010000;
            14'h6156: o_data_a = 16'b1110110010100000;
            14'h6157: o_data_a = 16'b1111000010001000;
            14'h6158: o_data_a = 16'b0000000000000011;
            14'h6159: o_data_a = 16'b1110110000010000;
            14'h615a: o_data_a = 16'b0000000000000000;
            14'h615b: o_data_a = 16'b1111110111101000;
            14'h615c: o_data_a = 16'b1110110010100000;
            14'h615d: o_data_a = 16'b1110001100001000;
            14'h615e: o_data_a = 16'b0000000000000000;
            14'h615f: o_data_a = 16'b1111110010101000;
            14'h6160: o_data_a = 16'b1111110000010000;
            14'h6161: o_data_a = 16'b1110110010100000;
            14'h6162: o_data_a = 16'b1111000010001000;
            14'h6163: o_data_a = 16'b0000000000000000;
            14'h6164: o_data_a = 16'b1111110010101000;
            14'h6165: o_data_a = 16'b1111110000010000;
            14'h6166: o_data_a = 16'b0000000000000001;
            14'h6167: o_data_a = 16'b1111110111100000;
            14'h6168: o_data_a = 16'b1110110111100000;
            14'h6169: o_data_a = 16'b1110001100001000;
            14'h616a: o_data_a = 16'b0110000111000110;
            14'h616b: o_data_a = 16'b1110101010000111;
            14'h616c: o_data_a = 16'b0000000000000001;
            14'h616d: o_data_a = 16'b1111110111100000;
            14'h616e: o_data_a = 16'b1110110111100000;
            14'h616f: o_data_a = 16'b1111110000010000;
            14'h6170: o_data_a = 16'b0000000000000000;
            14'h6171: o_data_a = 16'b1111110111101000;
            14'h6172: o_data_a = 16'b1110110010100000;
            14'h6173: o_data_a = 16'b1110001100001000;
            14'h6174: o_data_a = 16'b0000000000000010;
            14'h6175: o_data_a = 16'b1110110000010000;
            14'h6176: o_data_a = 16'b0000000000000000;
            14'h6177: o_data_a = 16'b1111110111101000;
            14'h6178: o_data_a = 16'b1110110010100000;
            14'h6179: o_data_a = 16'b1110001100001000;
            14'h617a: o_data_a = 16'b0000000000000001;
            14'h617b: o_data_a = 16'b1111110000100000;
            14'h617c: o_data_a = 16'b1111110000010000;
            14'h617d: o_data_a = 16'b0000000000000000;
            14'h617e: o_data_a = 16'b1111110111101000;
            14'h617f: o_data_a = 16'b1110110010100000;
            14'h6180: o_data_a = 16'b1110001100001000;
            14'h6181: o_data_a = 16'b0000000000000001;
            14'h6182: o_data_a = 16'b1111110111100000;
            14'h6183: o_data_a = 16'b1111110000010000;
            14'h6184: o_data_a = 16'b0000000000000000;
            14'h6185: o_data_a = 16'b1111110111101000;
            14'h6186: o_data_a = 16'b1110110010100000;
            14'h6187: o_data_a = 16'b1110001100001000;
            14'h6188: o_data_a = 16'b0000000000000000;
            14'h6189: o_data_a = 16'b1111110010101000;
            14'h618a: o_data_a = 16'b1111110000010000;
            14'h618b: o_data_a = 16'b1110110010100000;
            14'h618c: o_data_a = 16'b1111000111001000;
            14'h618d: o_data_a = 16'b0000000000000010;
            14'h618e: o_data_a = 16'b1110110000010000;
            14'h618f: o_data_a = 16'b0000000000001101;
            14'h6190: o_data_a = 16'b1110001100001000;
            14'h6191: o_data_a = 16'b0001101010100110;
            14'h6192: o_data_a = 16'b1110110000010000;
            14'h6193: o_data_a = 16'b0000000000001110;
            14'h6194: o_data_a = 16'b1110001100001000;
            14'h6195: o_data_a = 16'b0110000110011001;
            14'h6196: o_data_a = 16'b1110110000010000;
            14'h6197: o_data_a = 16'b0000000001011111;
            14'h6198: o_data_a = 16'b1110101010000111;
            14'h6199: o_data_a = 16'b0000000000000000;
            14'h619a: o_data_a = 16'b1111110010101000;
            14'h619b: o_data_a = 16'b1111110000010000;
            14'h619c: o_data_a = 16'b1110110010100000;
            14'h619d: o_data_a = 16'b1111000010001000;
            14'h619e: o_data_a = 16'b0000000000000101;
            14'h619f: o_data_a = 16'b1110110000010000;
            14'h61a0: o_data_a = 16'b0000000000000000;
            14'h61a1: o_data_a = 16'b1111110111101000;
            14'h61a2: o_data_a = 16'b1110110010100000;
            14'h61a3: o_data_a = 16'b1110001100001000;
            14'h61a4: o_data_a = 16'b0000000000000000;
            14'h61a5: o_data_a = 16'b1111110010101000;
            14'h61a6: o_data_a = 16'b1111110000010000;
            14'h61a7: o_data_a = 16'b1110110010100000;
            14'h61a8: o_data_a = 16'b1111000010001000;
            14'h61a9: o_data_a = 16'b0000000000000000;
            14'h61aa: o_data_a = 16'b1111110010101000;
            14'h61ab: o_data_a = 16'b1111110000010000;
            14'h61ac: o_data_a = 16'b0000000000000001;
            14'h61ad: o_data_a = 16'b1111110111100000;
            14'h61ae: o_data_a = 16'b1110110111100000;
            14'h61af: o_data_a = 16'b1110001100001000;
            14'h61b0: o_data_a = 16'b0000000000000001;
            14'h61b1: o_data_a = 16'b1111110111100000;
            14'h61b2: o_data_a = 16'b1111110000010000;
            14'h61b3: o_data_a = 16'b0000000000000000;
            14'h61b4: o_data_a = 16'b1111110111101000;
            14'h61b5: o_data_a = 16'b1110110010100000;
            14'h61b6: o_data_a = 16'b1110001100001000;
            14'h61b7: o_data_a = 16'b0000000000000000;
            14'h61b8: o_data_a = 16'b1111110111001000;
            14'h61b9: o_data_a = 16'b1111110010100000;
            14'h61ba: o_data_a = 16'b1110111111001000;
            14'h61bb: o_data_a = 16'b0000000000000000;
            14'h61bc: o_data_a = 16'b1111110010101000;
            14'h61bd: o_data_a = 16'b1111110000010000;
            14'h61be: o_data_a = 16'b1110110010100000;
            14'h61bf: o_data_a = 16'b1111000111001000;
            14'h61c0: o_data_a = 16'b0000000000000000;
            14'h61c1: o_data_a = 16'b1111110010101000;
            14'h61c2: o_data_a = 16'b1111110000010000;
            14'h61c3: o_data_a = 16'b0000000000000001;
            14'h61c4: o_data_a = 16'b1111110111100000;
            14'h61c5: o_data_a = 16'b1110001100001000;
            14'h61c6: o_data_a = 16'b0000000000000001;
            14'h61c7: o_data_a = 16'b1111110000100000;
            14'h61c8: o_data_a = 16'b1111110000010000;
            14'h61c9: o_data_a = 16'b0000000000000000;
            14'h61ca: o_data_a = 16'b1111110111101000;
            14'h61cb: o_data_a = 16'b1110110010100000;
            14'h61cc: o_data_a = 16'b1110001100001000;
            14'h61cd: o_data_a = 16'b0000000000000000;
            14'h61ce: o_data_a = 16'b1111110111001000;
            14'h61cf: o_data_a = 16'b1111110010100000;
            14'h61d0: o_data_a = 16'b1110111111001000;
            14'h61d1: o_data_a = 16'b0000000000000000;
            14'h61d2: o_data_a = 16'b1111110010101000;
            14'h61d3: o_data_a = 16'b1111110000010000;
            14'h61d4: o_data_a = 16'b1110110010100000;
            14'h61d5: o_data_a = 16'b1111000010001000;
            14'h61d6: o_data_a = 16'b0000000000000000;
            14'h61d7: o_data_a = 16'b1111110010101000;
            14'h61d8: o_data_a = 16'b1111110000010000;
            14'h61d9: o_data_a = 16'b0000000000000001;
            14'h61da: o_data_a = 16'b1111110000100000;
            14'h61db: o_data_a = 16'b1110001100001000;
            14'h61dc: o_data_a = 16'b0000000000000010;
            14'h61dd: o_data_a = 16'b1111110000100000;
            14'h61de: o_data_a = 16'b1111110000010000;
            14'h61df: o_data_a = 16'b0000000000000000;
            14'h61e0: o_data_a = 16'b1111110111101000;
            14'h61e1: o_data_a = 16'b1110110010100000;
            14'h61e2: o_data_a = 16'b1110001100001000;
            14'h61e3: o_data_a = 16'b0000000000000010;
            14'h61e4: o_data_a = 16'b1111110111100000;
            14'h61e5: o_data_a = 16'b1111110000010000;
            14'h61e6: o_data_a = 16'b0000000000000000;
            14'h61e7: o_data_a = 16'b1111110111101000;
            14'h61e8: o_data_a = 16'b1110110010100000;
            14'h61e9: o_data_a = 16'b1110001100001000;
            14'h61ea: o_data_a = 16'b0000000000000001;
            14'h61eb: o_data_a = 16'b1111110000100000;
            14'h61ec: o_data_a = 16'b1111110000010000;
            14'h61ed: o_data_a = 16'b0000000000000000;
            14'h61ee: o_data_a = 16'b1111110111101000;
            14'h61ef: o_data_a = 16'b1110110010100000;
            14'h61f0: o_data_a = 16'b1110001100001000;
            14'h61f1: o_data_a = 16'b0000000000000001;
            14'h61f2: o_data_a = 16'b1111110111100000;
            14'h61f3: o_data_a = 16'b1111110000010000;
            14'h61f4: o_data_a = 16'b0000000000000000;
            14'h61f5: o_data_a = 16'b1111110111101000;
            14'h61f6: o_data_a = 16'b1110110010100000;
            14'h61f7: o_data_a = 16'b1110001100001000;
            14'h61f8: o_data_a = 16'b0000000000000100;
            14'h61f9: o_data_a = 16'b1110110000010000;
            14'h61fa: o_data_a = 16'b0000000000001101;
            14'h61fb: o_data_a = 16'b1110001100001000;
            14'h61fc: o_data_a = 16'b0101111001010111;
            14'h61fd: o_data_a = 16'b1110110000010000;
            14'h61fe: o_data_a = 16'b0000000000001110;
            14'h61ff: o_data_a = 16'b1110001100001000;
            14'h6200: o_data_a = 16'b0110001000000100;
            14'h6201: o_data_a = 16'b1110110000010000;
            14'h6202: o_data_a = 16'b0000000001011111;
            14'h6203: o_data_a = 16'b1110101010000111;
            14'h6204: o_data_a = 16'b0000000000000000;
            14'h6205: o_data_a = 16'b1111110010101000;
            14'h6206: o_data_a = 16'b1111110000010000;
            14'h6207: o_data_a = 16'b0000000000000101;
            14'h6208: o_data_a = 16'b1110001100001000;
            14'h6209: o_data_a = 16'b0110000100000001;
            14'h620a: o_data_a = 16'b1110101010000111;
            14'h620b: o_data_a = 16'b0000000000000000;
            14'h620c: o_data_a = 16'b1111110111001000;
            14'h620d: o_data_a = 16'b1111110010100000;
            14'h620e: o_data_a = 16'b1110101010001000;
            14'h620f: o_data_a = 16'b0000000000110110;
            14'h6210: o_data_a = 16'b1110101010000111;
            14'h6211: o_data_a = 16'b0000000000000011;
            14'h6212: o_data_a = 16'b1110110000010000;
            14'h6213: o_data_a = 16'b0000000000000000;
            14'h6214: o_data_a = 16'b1111110111101000;
            14'h6215: o_data_a = 16'b1110110010100000;
            14'h6216: o_data_a = 16'b1110001100001000;
            14'h6217: o_data_a = 16'b0000000000000001;
            14'h6218: o_data_a = 16'b1110110000010000;
            14'h6219: o_data_a = 16'b0000000000001101;
            14'h621a: o_data_a = 16'b1110001100001000;
            14'h621b: o_data_a = 16'b0010000111000011;
            14'h621c: o_data_a = 16'b1110110000010000;
            14'h621d: o_data_a = 16'b0000000000001110;
            14'h621e: o_data_a = 16'b1110001100001000;
            14'h621f: o_data_a = 16'b0110001000100011;
            14'h6220: o_data_a = 16'b1110110000010000;
            14'h6221: o_data_a = 16'b0000000001011111;
            14'h6222: o_data_a = 16'b1110101010000111;
            14'h6223: o_data_a = 16'b0000000000000000;
            14'h6224: o_data_a = 16'b1111110010101000;
            14'h6225: o_data_a = 16'b1111110000010000;
            14'h6226: o_data_a = 16'b0000000000000011;
            14'h6227: o_data_a = 16'b1110001100001000;
            14'h6228: o_data_a = 16'b0000000000000010;
            14'h6229: o_data_a = 16'b1111110000100000;
            14'h622a: o_data_a = 16'b1111110000010000;
            14'h622b: o_data_a = 16'b0000000000000000;
            14'h622c: o_data_a = 16'b1111110111101000;
            14'h622d: o_data_a = 16'b1110110010100000;
            14'h622e: o_data_a = 16'b1110001100001000;
            14'h622f: o_data_a = 16'b0000000000000000;
            14'h6230: o_data_a = 16'b1111110111001000;
            14'h6231: o_data_a = 16'b1111110010100000;
            14'h6232: o_data_a = 16'b1110101010001000;
            14'h6233: o_data_a = 16'b0110001000110111;
            14'h6234: o_data_a = 16'b1110110000010000;
            14'h6235: o_data_a = 16'b0000000000100110;
            14'h6236: o_data_a = 16'b1110101010000111;
            14'h6237: o_data_a = 16'b0000000000000000;
            14'h6238: o_data_a = 16'b1111110010101000;
            14'h6239: o_data_a = 16'b1111110000010000;
            14'h623a: o_data_a = 16'b0110001000111110;
            14'h623b: o_data_a = 16'b1110001100000101;
            14'h623c: o_data_a = 16'b0110001001010101;
            14'h623d: o_data_a = 16'b1110101010000111;
            14'h623e: o_data_a = 16'b0000000000001110;
            14'h623f: o_data_a = 16'b1110110000010000;
            14'h6240: o_data_a = 16'b0000000000000000;
            14'h6241: o_data_a = 16'b1111110111101000;
            14'h6242: o_data_a = 16'b1110110010100000;
            14'h6243: o_data_a = 16'b1110001100001000;
            14'h6244: o_data_a = 16'b0000000000000001;
            14'h6245: o_data_a = 16'b1110110000010000;
            14'h6246: o_data_a = 16'b0000000000001101;
            14'h6247: o_data_a = 16'b1110001100001000;
            14'h6248: o_data_a = 16'b0110101011011001;
            14'h6249: o_data_a = 16'b1110110000010000;
            14'h624a: o_data_a = 16'b0000000000001110;
            14'h624b: o_data_a = 16'b1110001100001000;
            14'h624c: o_data_a = 16'b0110001001010000;
            14'h624d: o_data_a = 16'b1110110000010000;
            14'h624e: o_data_a = 16'b0000000001011111;
            14'h624f: o_data_a = 16'b1110101010000111;
            14'h6250: o_data_a = 16'b0000000000000000;
            14'h6251: o_data_a = 16'b1111110010101000;
            14'h6252: o_data_a = 16'b1111110000010000;
            14'h6253: o_data_a = 16'b0000000000000101;
            14'h6254: o_data_a = 16'b1110001100001000;
            14'h6255: o_data_a = 16'b0000000000000010;
            14'h6256: o_data_a = 16'b1111110000100000;
            14'h6257: o_data_a = 16'b1111110000010000;
            14'h6258: o_data_a = 16'b0000000000000000;
            14'h6259: o_data_a = 16'b1111110111101000;
            14'h625a: o_data_a = 16'b1110110010100000;
            14'h625b: o_data_a = 16'b1110001100001000;
            14'h625c: o_data_a = 16'b0000000000000000;
            14'h625d: o_data_a = 16'b1111110111001000;
            14'h625e: o_data_a = 16'b1111110010100000;
            14'h625f: o_data_a = 16'b1110101010001000;
            14'h6260: o_data_a = 16'b0110001001100100;
            14'h6261: o_data_a = 16'b1110110000010000;
            14'h6262: o_data_a = 16'b0000000000010110;
            14'h6263: o_data_a = 16'b1110101010000111;
            14'h6264: o_data_a = 16'b0000000000000000;
            14'h6265: o_data_a = 16'b1111110010101000;
            14'h6266: o_data_a = 16'b1111110000010000;
            14'h6267: o_data_a = 16'b0110001001101011;
            14'h6268: o_data_a = 16'b1110001100000101;
            14'h6269: o_data_a = 16'b0110001010000100;
            14'h626a: o_data_a = 16'b1110101010000111;
            14'h626b: o_data_a = 16'b0000000000000010;
            14'h626c: o_data_a = 16'b1111110000100000;
            14'h626d: o_data_a = 16'b1111110000010000;
            14'h626e: o_data_a = 16'b0000000000000000;
            14'h626f: o_data_a = 16'b1111110111101000;
            14'h6270: o_data_a = 16'b1110110010100000;
            14'h6271: o_data_a = 16'b1110001100001000;
            14'h6272: o_data_a = 16'b0000000000000001;
            14'h6273: o_data_a = 16'b1110110000010000;
            14'h6274: o_data_a = 16'b0000000000001101;
            14'h6275: o_data_a = 16'b1110001100001000;
            14'h6276: o_data_a = 16'b0001011010110000;
            14'h6277: o_data_a = 16'b1110110000010000;
            14'h6278: o_data_a = 16'b0000000000001110;
            14'h6279: o_data_a = 16'b1110001100001000;
            14'h627a: o_data_a = 16'b0110001001111110;
            14'h627b: o_data_a = 16'b1110110000010000;
            14'h627c: o_data_a = 16'b0000000001011111;
            14'h627d: o_data_a = 16'b1110101010000111;
            14'h627e: o_data_a = 16'b0000000000000000;
            14'h627f: o_data_a = 16'b1111110010101000;
            14'h6280: o_data_a = 16'b1111110000010000;
            14'h6281: o_data_a = 16'b0000000000000011;
            14'h6282: o_data_a = 16'b1111110111100000;
            14'h6283: o_data_a = 16'b1110001100001000;
            14'h6284: o_data_a = 16'b0000000000000010;
            14'h6285: o_data_a = 16'b1111110000100000;
            14'h6286: o_data_a = 16'b1111110000010000;
            14'h6287: o_data_a = 16'b0000000000000000;
            14'h6288: o_data_a = 16'b1111110111101000;
            14'h6289: o_data_a = 16'b1110110010100000;
            14'h628a: o_data_a = 16'b1110001100001000;
            14'h628b: o_data_a = 16'b0000000000000000;
            14'h628c: o_data_a = 16'b1111110010101000;
            14'h628d: o_data_a = 16'b1111110000010000;
            14'h628e: o_data_a = 16'b0000000000000011;
            14'h628f: o_data_a = 16'b1111110000100000;
            14'h6290: o_data_a = 16'b1110001100001000;
            14'h6291: o_data_a = 16'b0000000000000000;
            14'h6292: o_data_a = 16'b1111110111001000;
            14'h6293: o_data_a = 16'b1111110010100000;
            14'h6294: o_data_a = 16'b1110101010001000;
            14'h6295: o_data_a = 16'b0000000000000000;
            14'h6296: o_data_a = 16'b1111110010101000;
            14'h6297: o_data_a = 16'b1111110000010000;
            14'h6298: o_data_a = 16'b0000000000000011;
            14'h6299: o_data_a = 16'b1111110111100000;
            14'h629a: o_data_a = 16'b1110110111100000;
            14'h629b: o_data_a = 16'b1110001100001000;
            14'h629c: o_data_a = 16'b0000000000000011;
            14'h629d: o_data_a = 16'b1111110000010000;
            14'h629e: o_data_a = 16'b0000000000000000;
            14'h629f: o_data_a = 16'b1111110111101000;
            14'h62a0: o_data_a = 16'b1110110010100000;
            14'h62a1: o_data_a = 16'b1110001100001000;
            14'h62a2: o_data_a = 16'b0000000000110110;
            14'h62a3: o_data_a = 16'b1110101010000111;
            14'h62a4: o_data_a = 16'b0000000000000010;
            14'h62a5: o_data_a = 16'b1111110000100000;
            14'h62a6: o_data_a = 16'b1111110000010000;
            14'h62a7: o_data_a = 16'b0000000000000000;
            14'h62a8: o_data_a = 16'b1111110111101000;
            14'h62a9: o_data_a = 16'b1110110010100000;
            14'h62aa: o_data_a = 16'b1110001100001000;
            14'h62ab: o_data_a = 16'b0000000000000000;
            14'h62ac: o_data_a = 16'b1111110010101000;
            14'h62ad: o_data_a = 16'b1111110000010000;
            14'h62ae: o_data_a = 16'b0000000000000011;
            14'h62af: o_data_a = 16'b1110001100001000;
            14'h62b0: o_data_a = 16'b0000000000000011;
            14'h62b1: o_data_a = 16'b1111110000100000;
            14'h62b2: o_data_a = 16'b1111110000010000;
            14'h62b3: o_data_a = 16'b0000000000000000;
            14'h62b4: o_data_a = 16'b1111110111101000;
            14'h62b5: o_data_a = 16'b1110110010100000;
            14'h62b6: o_data_a = 16'b1110001100001000;
            14'h62b7: o_data_a = 16'b0000000000000000;
            14'h62b8: o_data_a = 16'b1111110111001000;
            14'h62b9: o_data_a = 16'b1111110010100000;
            14'h62ba: o_data_a = 16'b1110101010001000;
            14'h62bb: o_data_a = 16'b0110001010111111;
            14'h62bc: o_data_a = 16'b1110110000010000;
            14'h62bd: o_data_a = 16'b0000000000010110;
            14'h62be: o_data_a = 16'b1110101010000111;
            14'h62bf: o_data_a = 16'b0000000000000000;
            14'h62c0: o_data_a = 16'b1111110010101000;
            14'h62c1: o_data_a = 16'b1111110000010000;
            14'h62c2: o_data_a = 16'b0110001011000110;
            14'h62c3: o_data_a = 16'b1110001100000101;
            14'h62c4: o_data_a = 16'b0110001011011110;
            14'h62c5: o_data_a = 16'b1110101010000111;
            14'h62c6: o_data_a = 16'b0000000000000011;
            14'h62c7: o_data_a = 16'b1111110111100000;
            14'h62c8: o_data_a = 16'b1111110000010000;
            14'h62c9: o_data_a = 16'b0000000000000000;
            14'h62ca: o_data_a = 16'b1111110111101000;
            14'h62cb: o_data_a = 16'b1110110010100000;
            14'h62cc: o_data_a = 16'b1110001100001000;
            14'h62cd: o_data_a = 16'b0000000000000001;
            14'h62ce: o_data_a = 16'b1110110000010000;
            14'h62cf: o_data_a = 16'b0000000000001101;
            14'h62d0: o_data_a = 16'b1110001100001000;
            14'h62d1: o_data_a = 16'b0001011011110101;
            14'h62d2: o_data_a = 16'b1110110000010000;
            14'h62d3: o_data_a = 16'b0000000000001110;
            14'h62d4: o_data_a = 16'b1110001100001000;
            14'h62d5: o_data_a = 16'b0110001011011001;
            14'h62d6: o_data_a = 16'b1110110000010000;
            14'h62d7: o_data_a = 16'b0000000001011111;
            14'h62d8: o_data_a = 16'b1110101010000111;
            14'h62d9: o_data_a = 16'b0000000000000000;
            14'h62da: o_data_a = 16'b1111110010101000;
            14'h62db: o_data_a = 16'b1111110000010000;
            14'h62dc: o_data_a = 16'b0000000000000101;
            14'h62dd: o_data_a = 16'b1110001100001000;
            14'h62de: o_data_a = 16'b0000000000000011;
            14'h62df: o_data_a = 16'b1111110000010000;
            14'h62e0: o_data_a = 16'b0000000000000000;
            14'h62e1: o_data_a = 16'b1111110111101000;
            14'h62e2: o_data_a = 16'b1110110010100000;
            14'h62e3: o_data_a = 16'b1110001100001000;
            14'h62e4: o_data_a = 16'b0000000000000001;
            14'h62e5: o_data_a = 16'b1110110000010000;
            14'h62e6: o_data_a = 16'b0000000000001101;
            14'h62e7: o_data_a = 16'b1110001100001000;
            14'h62e8: o_data_a = 16'b0010010010001101;
            14'h62e9: o_data_a = 16'b1110110000010000;
            14'h62ea: o_data_a = 16'b0000000000001110;
            14'h62eb: o_data_a = 16'b1110001100001000;
            14'h62ec: o_data_a = 16'b0110001011110000;
            14'h62ed: o_data_a = 16'b1110110000010000;
            14'h62ee: o_data_a = 16'b0000000001011111;
            14'h62ef: o_data_a = 16'b1110101010000111;
            14'h62f0: o_data_a = 16'b0000000000000000;
            14'h62f1: o_data_a = 16'b1111110010101000;
            14'h62f2: o_data_a = 16'b1111110000010000;
            14'h62f3: o_data_a = 16'b0000000000000101;
            14'h62f4: o_data_a = 16'b1110001100001000;
            14'h62f5: o_data_a = 16'b0000000000000000;
            14'h62f6: o_data_a = 16'b1111110111001000;
            14'h62f7: o_data_a = 16'b1111110010100000;
            14'h62f8: o_data_a = 16'b1110101010001000;
            14'h62f9: o_data_a = 16'b0000000000110110;
            14'h62fa: o_data_a = 16'b1110101010000111;
            14'h62fb: o_data_a = 16'b0000000000000010;
            14'h62fc: o_data_a = 16'b1111110000100000;
            14'h62fd: o_data_a = 16'b1111110000010000;
            14'h62fe: o_data_a = 16'b0000000000000000;
            14'h62ff: o_data_a = 16'b1111110111101000;
            14'h6300: o_data_a = 16'b1110110010100000;
            14'h6301: o_data_a = 16'b1110001100001000;
            14'h6302: o_data_a = 16'b0000000000000000;
            14'h6303: o_data_a = 16'b1111110010101000;
            14'h6304: o_data_a = 16'b1111110000010000;
            14'h6305: o_data_a = 16'b0000000000000011;
            14'h6306: o_data_a = 16'b1110001100001000;
            14'h6307: o_data_a = 16'b0000000000000011;
            14'h6308: o_data_a = 16'b1111110111100000;
            14'h6309: o_data_a = 16'b1110110111100000;
            14'h630a: o_data_a = 16'b1111110000010000;
            14'h630b: o_data_a = 16'b0000000000000000;
            14'h630c: o_data_a = 16'b1111110111101000;
            14'h630d: o_data_a = 16'b1110110010100000;
            14'h630e: o_data_a = 16'b1110001100001000;
            14'h630f: o_data_a = 16'b0000000000110110;
            14'h6310: o_data_a = 16'b1110101010000111;
            14'h6311: o_data_a = 16'b0000000000000010;
            14'h6312: o_data_a = 16'b1111110000100000;
            14'h6313: o_data_a = 16'b1111110000010000;
            14'h6314: o_data_a = 16'b0000000000000000;
            14'h6315: o_data_a = 16'b1111110111101000;
            14'h6316: o_data_a = 16'b1110110010100000;
            14'h6317: o_data_a = 16'b1110001100001000;
            14'h6318: o_data_a = 16'b0000000000000000;
            14'h6319: o_data_a = 16'b1111110010101000;
            14'h631a: o_data_a = 16'b1111110000010000;
            14'h631b: o_data_a = 16'b0000000000000011;
            14'h631c: o_data_a = 16'b1110001100001000;
            14'h631d: o_data_a = 16'b0000000000000010;
            14'h631e: o_data_a = 16'b1111110111100000;
            14'h631f: o_data_a = 16'b1111110000010000;
            14'h6320: o_data_a = 16'b0000000000000000;
            14'h6321: o_data_a = 16'b1111110111101000;
            14'h6322: o_data_a = 16'b1110110010100000;
            14'h6323: o_data_a = 16'b1110001100001000;
            14'h6324: o_data_a = 16'b0000000000000000;
            14'h6325: o_data_a = 16'b1111110111001000;
            14'h6326: o_data_a = 16'b1111110010100000;
            14'h6327: o_data_a = 16'b1110101010001000;
            14'h6328: o_data_a = 16'b0110001100101100;
            14'h6329: o_data_a = 16'b1110110000010000;
            14'h632a: o_data_a = 16'b0000000000100110;
            14'h632b: o_data_a = 16'b1110101010000111;
            14'h632c: o_data_a = 16'b0000000000000010;
            14'h632d: o_data_a = 16'b1111110111100000;
            14'h632e: o_data_a = 16'b1111110000010000;
            14'h632f: o_data_a = 16'b0000000000000000;
            14'h6330: o_data_a = 16'b1111110111101000;
            14'h6331: o_data_a = 16'b1110110010100000;
            14'h6332: o_data_a = 16'b1110001100001000;
            14'h6333: o_data_a = 16'b0000000000000011;
            14'h6334: o_data_a = 16'b1111110111100000;
            14'h6335: o_data_a = 16'b1110110111100000;
            14'h6336: o_data_a = 16'b1111110000010000;
            14'h6337: o_data_a = 16'b0000000000000000;
            14'h6338: o_data_a = 16'b1111110111101000;
            14'h6339: o_data_a = 16'b1110110010100000;
            14'h633a: o_data_a = 16'b1110001100001000;
            14'h633b: o_data_a = 16'b0110001100111111;
            14'h633c: o_data_a = 16'b1110110000010000;
            14'h633d: o_data_a = 16'b0000000000010110;
            14'h633e: o_data_a = 16'b1110101010000111;
            14'h633f: o_data_a = 16'b0000000000000000;
            14'h6340: o_data_a = 16'b1111110010101000;
            14'h6341: o_data_a = 16'b1111110000010000;
            14'h6342: o_data_a = 16'b1110110010100000;
            14'h6343: o_data_a = 16'b1111010101001000;
            14'h6344: o_data_a = 16'b0000000000000010;
            14'h6345: o_data_a = 16'b1111110111100000;
            14'h6346: o_data_a = 16'b1111110000010000;
            14'h6347: o_data_a = 16'b0000000000000000;
            14'h6348: o_data_a = 16'b1111110111101000;
            14'h6349: o_data_a = 16'b1110110010100000;
            14'h634a: o_data_a = 16'b1110001100001000;
            14'h634b: o_data_a = 16'b0000000000000011;
            14'h634c: o_data_a = 16'b1111110111100000;
            14'h634d: o_data_a = 16'b1110110111100000;
            14'h634e: o_data_a = 16'b1111110000010000;
            14'h634f: o_data_a = 16'b0000000000000000;
            14'h6350: o_data_a = 16'b1111110111101000;
            14'h6351: o_data_a = 16'b1110110010100000;
            14'h6352: o_data_a = 16'b1110001100001000;
            14'h6353: o_data_a = 16'b0110001101010111;
            14'h6354: o_data_a = 16'b1110110000010000;
            14'h6355: o_data_a = 16'b0000000000000110;
            14'h6356: o_data_a = 16'b1110101010000111;
            14'h6357: o_data_a = 16'b0000000000000000;
            14'h6358: o_data_a = 16'b1111110010101000;
            14'h6359: o_data_a = 16'b1111110000010000;
            14'h635a: o_data_a = 16'b1110110010100000;
            14'h635b: o_data_a = 16'b1111010101001000;
            14'h635c: o_data_a = 16'b0000000000000000;
            14'h635d: o_data_a = 16'b1111110010101000;
            14'h635e: o_data_a = 16'b1111110000010000;
            14'h635f: o_data_a = 16'b0110001101100011;
            14'h6360: o_data_a = 16'b1110001100000101;
            14'h6361: o_data_a = 16'b0110001101111010;
            14'h6362: o_data_a = 16'b1110101010000111;
            14'h6363: o_data_a = 16'b0000000000001111;
            14'h6364: o_data_a = 16'b1110110000010000;
            14'h6365: o_data_a = 16'b0000000000000000;
            14'h6366: o_data_a = 16'b1111110111101000;
            14'h6367: o_data_a = 16'b1110110010100000;
            14'h6368: o_data_a = 16'b1110001100001000;
            14'h6369: o_data_a = 16'b0000000000000001;
            14'h636a: o_data_a = 16'b1110110000010000;
            14'h636b: o_data_a = 16'b0000000000001101;
            14'h636c: o_data_a = 16'b1110001100001000;
            14'h636d: o_data_a = 16'b0110101011011001;
            14'h636e: o_data_a = 16'b1110110000010000;
            14'h636f: o_data_a = 16'b0000000000001110;
            14'h6370: o_data_a = 16'b1110001100001000;
            14'h6371: o_data_a = 16'b0110001101110101;
            14'h6372: o_data_a = 16'b1110110000010000;
            14'h6373: o_data_a = 16'b0000000001011111;
            14'h6374: o_data_a = 16'b1110101010000111;
            14'h6375: o_data_a = 16'b0000000000000000;
            14'h6376: o_data_a = 16'b1111110010101000;
            14'h6377: o_data_a = 16'b1111110000010000;
            14'h6378: o_data_a = 16'b0000000000000101;
            14'h6379: o_data_a = 16'b1110001100001000;
            14'h637a: o_data_a = 16'b0000000000000010;
            14'h637b: o_data_a = 16'b1111110111100000;
            14'h637c: o_data_a = 16'b1111110000010000;
            14'h637d: o_data_a = 16'b0000000000000000;
            14'h637e: o_data_a = 16'b1111110111101000;
            14'h637f: o_data_a = 16'b1110110010100000;
            14'h6380: o_data_a = 16'b1110001100001000;
            14'h6381: o_data_a = 16'b0000000000000011;
            14'h6382: o_data_a = 16'b1111110111100000;
            14'h6383: o_data_a = 16'b1111110000010000;
            14'h6384: o_data_a = 16'b0000000000000000;
            14'h6385: o_data_a = 16'b1111110111101000;
            14'h6386: o_data_a = 16'b1110110010100000;
            14'h6387: o_data_a = 16'b1110001100001000;
            14'h6388: o_data_a = 16'b0000000000000000;
            14'h6389: o_data_a = 16'b1111110010101000;
            14'h638a: o_data_a = 16'b1111110000010000;
            14'h638b: o_data_a = 16'b1110110010100000;
            14'h638c: o_data_a = 16'b1111000010001000;
            14'h638d: o_data_a = 16'b0000000000000000;
            14'h638e: o_data_a = 16'b1111110010101000;
            14'h638f: o_data_a = 16'b1111110000010000;
            14'h6390: o_data_a = 16'b0000000000000100;
            14'h6391: o_data_a = 16'b1110001100001000;
            14'h6392: o_data_a = 16'b0000000000000100;
            14'h6393: o_data_a = 16'b1111110000100000;
            14'h6394: o_data_a = 16'b1111110000010000;
            14'h6395: o_data_a = 16'b0000000000000000;
            14'h6396: o_data_a = 16'b1111110111101000;
            14'h6397: o_data_a = 16'b1110110010100000;
            14'h6398: o_data_a = 16'b1110001100001000;
            14'h6399: o_data_a = 16'b0000000000110110;
            14'h639a: o_data_a = 16'b1110101010000111;
            14'h639b: o_data_a = 16'b0000000000000010;
            14'h639c: o_data_a = 16'b1111110000100000;
            14'h639d: o_data_a = 16'b1111110000010000;
            14'h639e: o_data_a = 16'b0000000000000000;
            14'h639f: o_data_a = 16'b1111110111101000;
            14'h63a0: o_data_a = 16'b1110110010100000;
            14'h63a1: o_data_a = 16'b1110001100001000;
            14'h63a2: o_data_a = 16'b0000000000000000;
            14'h63a3: o_data_a = 16'b1111110010101000;
            14'h63a4: o_data_a = 16'b1111110000010000;
            14'h63a5: o_data_a = 16'b0000000000000011;
            14'h63a6: o_data_a = 16'b1110001100001000;
            14'h63a7: o_data_a = 16'b0000000000000010;
            14'h63a8: o_data_a = 16'b1111110111100000;
            14'h63a9: o_data_a = 16'b1111110000010000;
            14'h63aa: o_data_a = 16'b0000000000000000;
            14'h63ab: o_data_a = 16'b1111110111101000;
            14'h63ac: o_data_a = 16'b1110110010100000;
            14'h63ad: o_data_a = 16'b1110001100001000;
            14'h63ae: o_data_a = 16'b0000000000000000;
            14'h63af: o_data_a = 16'b1111110111001000;
            14'h63b0: o_data_a = 16'b1111110010100000;
            14'h63b1: o_data_a = 16'b1110101010001000;
            14'h63b2: o_data_a = 16'b0110001110110110;
            14'h63b3: o_data_a = 16'b1110110000010000;
            14'h63b4: o_data_a = 16'b0000000000100110;
            14'h63b5: o_data_a = 16'b1110101010000111;
            14'h63b6: o_data_a = 16'b0000000000000010;
            14'h63b7: o_data_a = 16'b1111110111100000;
            14'h63b8: o_data_a = 16'b1111110000010000;
            14'h63b9: o_data_a = 16'b0000000000000000;
            14'h63ba: o_data_a = 16'b1111110111101000;
            14'h63bb: o_data_a = 16'b1110110010100000;
            14'h63bc: o_data_a = 16'b1110001100001000;
            14'h63bd: o_data_a = 16'b0000000000000011;
            14'h63be: o_data_a = 16'b1111110111100000;
            14'h63bf: o_data_a = 16'b1110110111100000;
            14'h63c0: o_data_a = 16'b1111110000010000;
            14'h63c1: o_data_a = 16'b0000000000000000;
            14'h63c2: o_data_a = 16'b1111110111101000;
            14'h63c3: o_data_a = 16'b1110110010100000;
            14'h63c4: o_data_a = 16'b1110001100001000;
            14'h63c5: o_data_a = 16'b0110001111001001;
            14'h63c6: o_data_a = 16'b1110110000010000;
            14'h63c7: o_data_a = 16'b0000000000010110;
            14'h63c8: o_data_a = 16'b1110101010000111;
            14'h63c9: o_data_a = 16'b0000000000000000;
            14'h63ca: o_data_a = 16'b1111110010101000;
            14'h63cb: o_data_a = 16'b1111110000010000;
            14'h63cc: o_data_a = 16'b1110110010100000;
            14'h63cd: o_data_a = 16'b1111010101001000;
            14'h63ce: o_data_a = 16'b0000000000000010;
            14'h63cf: o_data_a = 16'b1111110111100000;
            14'h63d0: o_data_a = 16'b1111110000010000;
            14'h63d1: o_data_a = 16'b0000000000000000;
            14'h63d2: o_data_a = 16'b1111110111101000;
            14'h63d3: o_data_a = 16'b1110110010100000;
            14'h63d4: o_data_a = 16'b1110001100001000;
            14'h63d5: o_data_a = 16'b0000000000000011;
            14'h63d6: o_data_a = 16'b1111110111100000;
            14'h63d7: o_data_a = 16'b1110110111100000;
            14'h63d8: o_data_a = 16'b1111110000010000;
            14'h63d9: o_data_a = 16'b0000000000000000;
            14'h63da: o_data_a = 16'b1111110111101000;
            14'h63db: o_data_a = 16'b1110110010100000;
            14'h63dc: o_data_a = 16'b1110001100001000;
            14'h63dd: o_data_a = 16'b0110001111100001;
            14'h63de: o_data_a = 16'b1110110000010000;
            14'h63df: o_data_a = 16'b0000000000000110;
            14'h63e0: o_data_a = 16'b1110101010000111;
            14'h63e1: o_data_a = 16'b0000000000000000;
            14'h63e2: o_data_a = 16'b1111110010101000;
            14'h63e3: o_data_a = 16'b1111110000010000;
            14'h63e4: o_data_a = 16'b1110110010100000;
            14'h63e5: o_data_a = 16'b1111010101001000;
            14'h63e6: o_data_a = 16'b0000000000000000;
            14'h63e7: o_data_a = 16'b1111110010101000;
            14'h63e8: o_data_a = 16'b1111110000010000;
            14'h63e9: o_data_a = 16'b0110001111101101;
            14'h63ea: o_data_a = 16'b1110001100000101;
            14'h63eb: o_data_a = 16'b0110010000000100;
            14'h63ec: o_data_a = 16'b1110101010000111;
            14'h63ed: o_data_a = 16'b0000000000010000;
            14'h63ee: o_data_a = 16'b1110110000010000;
            14'h63ef: o_data_a = 16'b0000000000000000;
            14'h63f0: o_data_a = 16'b1111110111101000;
            14'h63f1: o_data_a = 16'b1110110010100000;
            14'h63f2: o_data_a = 16'b1110001100001000;
            14'h63f3: o_data_a = 16'b0000000000000001;
            14'h63f4: o_data_a = 16'b1110110000010000;
            14'h63f5: o_data_a = 16'b0000000000001101;
            14'h63f6: o_data_a = 16'b1110001100001000;
            14'h63f7: o_data_a = 16'b0110101011011001;
            14'h63f8: o_data_a = 16'b1110110000010000;
            14'h63f9: o_data_a = 16'b0000000000001110;
            14'h63fa: o_data_a = 16'b1110001100001000;
            14'h63fb: o_data_a = 16'b0110001111111111;
            14'h63fc: o_data_a = 16'b1110110000010000;
            14'h63fd: o_data_a = 16'b0000000001011111;
            14'h63fe: o_data_a = 16'b1110101010000111;
            14'h63ff: o_data_a = 16'b0000000000000000;
            14'h6400: o_data_a = 16'b1111110010101000;
            14'h6401: o_data_a = 16'b1111110000010000;
            14'h6402: o_data_a = 16'b0000000000000101;
            14'h6403: o_data_a = 16'b1110001100001000;
            14'h6404: o_data_a = 16'b0000000000000010;
            14'h6405: o_data_a = 16'b1111110111100000;
            14'h6406: o_data_a = 16'b1111110000010000;
            14'h6407: o_data_a = 16'b0000000000000000;
            14'h6408: o_data_a = 16'b1111110111101000;
            14'h6409: o_data_a = 16'b1110110010100000;
            14'h640a: o_data_a = 16'b1110001100001000;
            14'h640b: o_data_a = 16'b0000000000000011;
            14'h640c: o_data_a = 16'b1111110111100000;
            14'h640d: o_data_a = 16'b1111110000010000;
            14'h640e: o_data_a = 16'b0000000000000000;
            14'h640f: o_data_a = 16'b1111110111101000;
            14'h6410: o_data_a = 16'b1110110010100000;
            14'h6411: o_data_a = 16'b1110001100001000;
            14'h6412: o_data_a = 16'b0000000000000000;
            14'h6413: o_data_a = 16'b1111110010101000;
            14'h6414: o_data_a = 16'b1111110000010000;
            14'h6415: o_data_a = 16'b1110110010100000;
            14'h6416: o_data_a = 16'b1111000010001000;
            14'h6417: o_data_a = 16'b0000000000000010;
            14'h6418: o_data_a = 16'b1111110111100000;
            14'h6419: o_data_a = 16'b1110110111100000;
            14'h641a: o_data_a = 16'b1111110000010000;
            14'h641b: o_data_a = 16'b0000000000000000;
            14'h641c: o_data_a = 16'b1111110111101000;
            14'h641d: o_data_a = 16'b1110110010100000;
            14'h641e: o_data_a = 16'b1110001100001000;
            14'h641f: o_data_a = 16'b0000000000000000;
            14'h6420: o_data_a = 16'b1111110010101000;
            14'h6421: o_data_a = 16'b1111110000010000;
            14'h6422: o_data_a = 16'b0000000000000101;
            14'h6423: o_data_a = 16'b1110001100001000;
            14'h6424: o_data_a = 16'b0000000000000000;
            14'h6425: o_data_a = 16'b1111110010101000;
            14'h6426: o_data_a = 16'b1111110000010000;
            14'h6427: o_data_a = 16'b0000000000000100;
            14'h6428: o_data_a = 16'b1110001100001000;
            14'h6429: o_data_a = 16'b0000000000000101;
            14'h642a: o_data_a = 16'b1111110000010000;
            14'h642b: o_data_a = 16'b0000000000000000;
            14'h642c: o_data_a = 16'b1111110111101000;
            14'h642d: o_data_a = 16'b1110110010100000;
            14'h642e: o_data_a = 16'b1110001100001000;
            14'h642f: o_data_a = 16'b0000000000000000;
            14'h6430: o_data_a = 16'b1111110010101000;
            14'h6431: o_data_a = 16'b1111110000010000;
            14'h6432: o_data_a = 16'b0000000000000100;
            14'h6433: o_data_a = 16'b1111110000100000;
            14'h6434: o_data_a = 16'b1110001100001000;
            14'h6435: o_data_a = 16'b0000000000000000;
            14'h6436: o_data_a = 16'b1111110111001000;
            14'h6437: o_data_a = 16'b1111110010100000;
            14'h6438: o_data_a = 16'b1110101010001000;
            14'h6439: o_data_a = 16'b0000000000110110;
            14'h643a: o_data_a = 16'b1110101010000111;
            14'h643b: o_data_a = 16'b0000000000000010;
            14'h643c: o_data_a = 16'b1111110000100000;
            14'h643d: o_data_a = 16'b1111110000010000;
            14'h643e: o_data_a = 16'b0000000000000000;
            14'h643f: o_data_a = 16'b1111110111101000;
            14'h6440: o_data_a = 16'b1110110010100000;
            14'h6441: o_data_a = 16'b1110001100001000;
            14'h6442: o_data_a = 16'b0000000000000000;
            14'h6443: o_data_a = 16'b1111110010101000;
            14'h6444: o_data_a = 16'b1111110000010000;
            14'h6445: o_data_a = 16'b0000000000000011;
            14'h6446: o_data_a = 16'b1110001100001000;
            14'h6447: o_data_a = 16'b0000000000000011;
            14'h6448: o_data_a = 16'b1111110111100000;
            14'h6449: o_data_a = 16'b1110110111100000;
            14'h644a: o_data_a = 16'b1111110000010000;
            14'h644b: o_data_a = 16'b0000000000000000;
            14'h644c: o_data_a = 16'b1111110111101000;
            14'h644d: o_data_a = 16'b1110110010100000;
            14'h644e: o_data_a = 16'b1110001100001000;
            14'h644f: o_data_a = 16'b0000000000000011;
            14'h6450: o_data_a = 16'b1111110000100000;
            14'h6451: o_data_a = 16'b1111110000010000;
            14'h6452: o_data_a = 16'b0000000000000000;
            14'h6453: o_data_a = 16'b1111110111101000;
            14'h6454: o_data_a = 16'b1110110010100000;
            14'h6455: o_data_a = 16'b1110001100001000;
            14'h6456: o_data_a = 16'b0110010001011010;
            14'h6457: o_data_a = 16'b1110110000010000;
            14'h6458: o_data_a = 16'b0000000000000110;
            14'h6459: o_data_a = 16'b1110101010000111;
            14'h645a: o_data_a = 16'b0000000000000000;
            14'h645b: o_data_a = 16'b1111110010101000;
            14'h645c: o_data_a = 16'b1111110000010000;
            14'h645d: o_data_a = 16'b0110010001100001;
            14'h645e: o_data_a = 16'b1110001100000101;
            14'h645f: o_data_a = 16'b0110010001111000;
            14'h6460: o_data_a = 16'b1110101010000111;
            14'h6461: o_data_a = 16'b0000000000010001;
            14'h6462: o_data_a = 16'b1110110000010000;
            14'h6463: o_data_a = 16'b0000000000000000;
            14'h6464: o_data_a = 16'b1111110111101000;
            14'h6465: o_data_a = 16'b1110110010100000;
            14'h6466: o_data_a = 16'b1110001100001000;
            14'h6467: o_data_a = 16'b0000000000000001;
            14'h6468: o_data_a = 16'b1110110000010000;
            14'h6469: o_data_a = 16'b0000000000001101;
            14'h646a: o_data_a = 16'b1110001100001000;
            14'h646b: o_data_a = 16'b0110101011011001;
            14'h646c: o_data_a = 16'b1110110000010000;
            14'h646d: o_data_a = 16'b0000000000001110;
            14'h646e: o_data_a = 16'b1110001100001000;
            14'h646f: o_data_a = 16'b0110010001110011;
            14'h6470: o_data_a = 16'b1110110000010000;
            14'h6471: o_data_a = 16'b0000000001011111;
            14'h6472: o_data_a = 16'b1110101010000111;
            14'h6473: o_data_a = 16'b0000000000000000;
            14'h6474: o_data_a = 16'b1111110010101000;
            14'h6475: o_data_a = 16'b1111110000010000;
            14'h6476: o_data_a = 16'b0000000000000101;
            14'h6477: o_data_a = 16'b1110001100001000;
            14'h6478: o_data_a = 16'b0000000000000011;
            14'h6479: o_data_a = 16'b1111110111100000;
            14'h647a: o_data_a = 16'b1110110111100000;
            14'h647b: o_data_a = 16'b1111110000010000;
            14'h647c: o_data_a = 16'b0000000000000000;
            14'h647d: o_data_a = 16'b1111110111101000;
            14'h647e: o_data_a = 16'b1110110010100000;
            14'h647f: o_data_a = 16'b1110001100001000;
            14'h6480: o_data_a = 16'b0000000000000011;
            14'h6481: o_data_a = 16'b1111110111100000;
            14'h6482: o_data_a = 16'b1111110000010000;
            14'h6483: o_data_a = 16'b0000000000000000;
            14'h6484: o_data_a = 16'b1111110111101000;
            14'h6485: o_data_a = 16'b1110110010100000;
            14'h6486: o_data_a = 16'b1110001100001000;
            14'h6487: o_data_a = 16'b0000000000000000;
            14'h6488: o_data_a = 16'b1111110010101000;
            14'h6489: o_data_a = 16'b1111110000010000;
            14'h648a: o_data_a = 16'b1110110010100000;
            14'h648b: o_data_a = 16'b1111000010001000;
            14'h648c: o_data_a = 16'b0000000000000010;
            14'h648d: o_data_a = 16'b1111110111100000;
            14'h648e: o_data_a = 16'b1111110000010000;
            14'h648f: o_data_a = 16'b0000000000000000;
            14'h6490: o_data_a = 16'b1111110111101000;
            14'h6491: o_data_a = 16'b1110110010100000;
            14'h6492: o_data_a = 16'b1110001100001000;
            14'h6493: o_data_a = 16'b0000000000000000;
            14'h6494: o_data_a = 16'b1111110010101000;
            14'h6495: o_data_a = 16'b1111110000010000;
            14'h6496: o_data_a = 16'b0000000000000101;
            14'h6497: o_data_a = 16'b1110001100001000;
            14'h6498: o_data_a = 16'b0000000000000000;
            14'h6499: o_data_a = 16'b1111110010101000;
            14'h649a: o_data_a = 16'b1111110000010000;
            14'h649b: o_data_a = 16'b0000000000000100;
            14'h649c: o_data_a = 16'b1110001100001000;
            14'h649d: o_data_a = 16'b0000000000000101;
            14'h649e: o_data_a = 16'b1111110000010000;
            14'h649f: o_data_a = 16'b0000000000000000;
            14'h64a0: o_data_a = 16'b1111110111101000;
            14'h64a1: o_data_a = 16'b1110110010100000;
            14'h64a2: o_data_a = 16'b1110001100001000;
            14'h64a3: o_data_a = 16'b0000000000000000;
            14'h64a4: o_data_a = 16'b1111110010101000;
            14'h64a5: o_data_a = 16'b1111110000010000;
            14'h64a6: o_data_a = 16'b0000000000000100;
            14'h64a7: o_data_a = 16'b1111110000100000;
            14'h64a8: o_data_a = 16'b1110001100001000;
            14'h64a9: o_data_a = 16'b0000000000000011;
            14'h64aa: o_data_a = 16'b1111110111100000;
            14'h64ab: o_data_a = 16'b1110110111100000;
            14'h64ac: o_data_a = 16'b1111110000010000;
            14'h64ad: o_data_a = 16'b0000000000000000;
            14'h64ae: o_data_a = 16'b1111110111101000;
            14'h64af: o_data_a = 16'b1110110010100000;
            14'h64b0: o_data_a = 16'b1110001100001000;
            14'h64b1: o_data_a = 16'b0000000000000000;
            14'h64b2: o_data_a = 16'b1111110111001000;
            14'h64b3: o_data_a = 16'b1111110010100000;
            14'h64b4: o_data_a = 16'b1110111111001000;
            14'h64b5: o_data_a = 16'b0000000000000000;
            14'h64b6: o_data_a = 16'b1111110010101000;
            14'h64b7: o_data_a = 16'b1111110000010000;
            14'h64b8: o_data_a = 16'b1110110010100000;
            14'h64b9: o_data_a = 16'b1111000010001000;
            14'h64ba: o_data_a = 16'b0000000000000000;
            14'h64bb: o_data_a = 16'b1111110010101000;
            14'h64bc: o_data_a = 16'b1111110000010000;
            14'h64bd: o_data_a = 16'b0000000000000011;
            14'h64be: o_data_a = 16'b1111110111100000;
            14'h64bf: o_data_a = 16'b1110110111100000;
            14'h64c0: o_data_a = 16'b1110001100001000;
            14'h64c1: o_data_a = 16'b0000000000000011;
            14'h64c2: o_data_a = 16'b1111110000010000;
            14'h64c3: o_data_a = 16'b0000000000000000;
            14'h64c4: o_data_a = 16'b1111110111101000;
            14'h64c5: o_data_a = 16'b1110110010100000;
            14'h64c6: o_data_a = 16'b1110001100001000;
            14'h64c7: o_data_a = 16'b0000000000110110;
            14'h64c8: o_data_a = 16'b1110101010000111;
            14'h64c9: o_data_a = 16'b0000000000000010;
            14'h64ca: o_data_a = 16'b1111110000100000;
            14'h64cb: o_data_a = 16'b1111110000010000;
            14'h64cc: o_data_a = 16'b0000000000000000;
            14'h64cd: o_data_a = 16'b1111110111101000;
            14'h64ce: o_data_a = 16'b1110110010100000;
            14'h64cf: o_data_a = 16'b1110001100001000;
            14'h64d0: o_data_a = 16'b0000000000000000;
            14'h64d1: o_data_a = 16'b1111110010101000;
            14'h64d2: o_data_a = 16'b1111110000010000;
            14'h64d3: o_data_a = 16'b0000000000000011;
            14'h64d4: o_data_a = 16'b1110001100001000;
            14'h64d5: o_data_a = 16'b0000000000000011;
            14'h64d6: o_data_a = 16'b1111110111100000;
            14'h64d7: o_data_a = 16'b1110110111100000;
            14'h64d8: o_data_a = 16'b1111110000010000;
            14'h64d9: o_data_a = 16'b0000000000000000;
            14'h64da: o_data_a = 16'b1111110111101000;
            14'h64db: o_data_a = 16'b1110110010100000;
            14'h64dc: o_data_a = 16'b1110001100001000;
            14'h64dd: o_data_a = 16'b0000000000000000;
            14'h64de: o_data_a = 16'b1111110111001000;
            14'h64df: o_data_a = 16'b1111110010100000;
            14'h64e0: o_data_a = 16'b1110101010001000;
            14'h64e1: o_data_a = 16'b0110010011100101;
            14'h64e2: o_data_a = 16'b1110110000010000;
            14'h64e3: o_data_a = 16'b0000000000000110;
            14'h64e4: o_data_a = 16'b1110101010000111;
            14'h64e5: o_data_a = 16'b0000000000000000;
            14'h64e6: o_data_a = 16'b1111110010101000;
            14'h64e7: o_data_a = 16'b1111110000010000;
            14'h64e8: o_data_a = 16'b0110010011101100;
            14'h64e9: o_data_a = 16'b1110001100000101;
            14'h64ea: o_data_a = 16'b0110010100000011;
            14'h64eb: o_data_a = 16'b1110101010000111;
            14'h64ec: o_data_a = 16'b0000000000010010;
            14'h64ed: o_data_a = 16'b1110110000010000;
            14'h64ee: o_data_a = 16'b0000000000000000;
            14'h64ef: o_data_a = 16'b1111110111101000;
            14'h64f0: o_data_a = 16'b1110110010100000;
            14'h64f1: o_data_a = 16'b1110001100001000;
            14'h64f2: o_data_a = 16'b0000000000000001;
            14'h64f3: o_data_a = 16'b1110110000010000;
            14'h64f4: o_data_a = 16'b0000000000001101;
            14'h64f5: o_data_a = 16'b1110001100001000;
            14'h64f6: o_data_a = 16'b0110101011011001;
            14'h64f7: o_data_a = 16'b1110110000010000;
            14'h64f8: o_data_a = 16'b0000000000001110;
            14'h64f9: o_data_a = 16'b1110001100001000;
            14'h64fa: o_data_a = 16'b0110010011111110;
            14'h64fb: o_data_a = 16'b1110110000010000;
            14'h64fc: o_data_a = 16'b0000000001011111;
            14'h64fd: o_data_a = 16'b1110101010000111;
            14'h64fe: o_data_a = 16'b0000000000000000;
            14'h64ff: o_data_a = 16'b1111110010101000;
            14'h6500: o_data_a = 16'b1111110000010000;
            14'h6501: o_data_a = 16'b0000000000000101;
            14'h6502: o_data_a = 16'b1110001100001000;
            14'h6503: o_data_a = 16'b0000000000000011;
            14'h6504: o_data_a = 16'b1111110111100000;
            14'h6505: o_data_a = 16'b1110110111100000;
            14'h6506: o_data_a = 16'b1111110000010000;
            14'h6507: o_data_a = 16'b0000000000000000;
            14'h6508: o_data_a = 16'b1111110111101000;
            14'h6509: o_data_a = 16'b1110110010100000;
            14'h650a: o_data_a = 16'b1110001100001000;
            14'h650b: o_data_a = 16'b0000000000000000;
            14'h650c: o_data_a = 16'b1111110111001000;
            14'h650d: o_data_a = 16'b1111110010100000;
            14'h650e: o_data_a = 16'b1110111111001000;
            14'h650f: o_data_a = 16'b0000000000000000;
            14'h6510: o_data_a = 16'b1111110010101000;
            14'h6511: o_data_a = 16'b1111110000010000;
            14'h6512: o_data_a = 16'b1110110010100000;
            14'h6513: o_data_a = 16'b1111000111001000;
            14'h6514: o_data_a = 16'b0000000000000000;
            14'h6515: o_data_a = 16'b1111110010101000;
            14'h6516: o_data_a = 16'b1111110000010000;
            14'h6517: o_data_a = 16'b0000000000000011;
            14'h6518: o_data_a = 16'b1111110111100000;
            14'h6519: o_data_a = 16'b1110110111100000;
            14'h651a: o_data_a = 16'b1110001100001000;
            14'h651b: o_data_a = 16'b0000000000000000;
            14'h651c: o_data_a = 16'b1111110111001000;
            14'h651d: o_data_a = 16'b1111110010100000;
            14'h651e: o_data_a = 16'b1110101010001000;
            14'h651f: o_data_a = 16'b0000000000110110;
            14'h6520: o_data_a = 16'b1110101010000111;
            14'h6521: o_data_a = 16'b0000000000000101;
            14'h6522: o_data_a = 16'b1110110000010000;
            14'h6523: o_data_a = 16'b1110001110010000;
            14'h6524: o_data_a = 16'b0000000000000000;
            14'h6525: o_data_a = 16'b1111110111101000;
            14'h6526: o_data_a = 16'b1110110010100000;
            14'h6527: o_data_a = 16'b1110101010001000;
            14'h6528: o_data_a = 16'b0110010100100011;
            14'h6529: o_data_a = 16'b1110001100000001;
            14'h652a: o_data_a = 16'b0000000000000010;
            14'h652b: o_data_a = 16'b1111110000100000;
            14'h652c: o_data_a = 16'b1111110000010000;
            14'h652d: o_data_a = 16'b0000000000000000;
            14'h652e: o_data_a = 16'b1111110111101000;
            14'h652f: o_data_a = 16'b1110110010100000;
            14'h6530: o_data_a = 16'b1110001100001000;
            14'h6531: o_data_a = 16'b0000000000000000;
            14'h6532: o_data_a = 16'b1111110010101000;
            14'h6533: o_data_a = 16'b1111110000010000;
            14'h6534: o_data_a = 16'b0000000000000011;
            14'h6535: o_data_a = 16'b1110001100001000;
            14'h6536: o_data_a = 16'b0000000000000011;
            14'h6537: o_data_a = 16'b1111110111100000;
            14'h6538: o_data_a = 16'b1110110111100000;
            14'h6539: o_data_a = 16'b1111110000010000;
            14'h653a: o_data_a = 16'b0000000000000000;
            14'h653b: o_data_a = 16'b1111110111101000;
            14'h653c: o_data_a = 16'b1110110010100000;
            14'h653d: o_data_a = 16'b1110001100001000;
            14'h653e: o_data_a = 16'b0000000000000000;
            14'h653f: o_data_a = 16'b1111110111001000;
            14'h6540: o_data_a = 16'b1111110010100000;
            14'h6541: o_data_a = 16'b1110101010001000;
            14'h6542: o_data_a = 16'b0110010101000110;
            14'h6543: o_data_a = 16'b1110110000010000;
            14'h6544: o_data_a = 16'b0000000000000110;
            14'h6545: o_data_a = 16'b1110101010000111;
            14'h6546: o_data_a = 16'b0000000000000000;
            14'h6547: o_data_a = 16'b1111110010101000;
            14'h6548: o_data_a = 16'b1111110000010000;
            14'h6549: o_data_a = 16'b0110010101001101;
            14'h654a: o_data_a = 16'b1110001100000101;
            14'h654b: o_data_a = 16'b0110010101010011;
            14'h654c: o_data_a = 16'b1110101010000111;
            14'h654d: o_data_a = 16'b0000000000000000;
            14'h654e: o_data_a = 16'b1111110111001000;
            14'h654f: o_data_a = 16'b1111110010100000;
            14'h6550: o_data_a = 16'b1110101010001000;
            14'h6551: o_data_a = 16'b0000000000110110;
            14'h6552: o_data_a = 16'b1110101010000111;
            14'h6553: o_data_a = 16'b0000000000000000;
            14'h6554: o_data_a = 16'b1111110111001000;
            14'h6555: o_data_a = 16'b1111110010100000;
            14'h6556: o_data_a = 16'b1110101010001000;
            14'h6557: o_data_a = 16'b0000000000000000;
            14'h6558: o_data_a = 16'b1111110010100000;
            14'h6559: o_data_a = 16'b1111110001001000;
            14'h655a: o_data_a = 16'b0000000000000000;
            14'h655b: o_data_a = 16'b1111110010101000;
            14'h655c: o_data_a = 16'b1111110000010000;
            14'h655d: o_data_a = 16'b0000000000000001;
            14'h655e: o_data_a = 16'b1111110111100000;
            14'h655f: o_data_a = 16'b1110110111100000;
            14'h6560: o_data_a = 16'b1110110111100000;
            14'h6561: o_data_a = 16'b1110001100001000;
            14'h6562: o_data_a = 16'b0000000000000000;
            14'h6563: o_data_a = 16'b1111110111001000;
            14'h6564: o_data_a = 16'b1111110010100000;
            14'h6565: o_data_a = 16'b1110101010001000;
            14'h6566: o_data_a = 16'b0000000000000011;
            14'h6567: o_data_a = 16'b1111110111100000;
            14'h6568: o_data_a = 16'b1111110000010000;
            14'h6569: o_data_a = 16'b0000000000000000;
            14'h656a: o_data_a = 16'b1111110111101000;
            14'h656b: o_data_a = 16'b1110110010100000;
            14'h656c: o_data_a = 16'b1110001100001000;
            14'h656d: o_data_a = 16'b0000000000000000;
            14'h656e: o_data_a = 16'b1111110010101000;
            14'h656f: o_data_a = 16'b1111110000010000;
            14'h6570: o_data_a = 16'b1110110010100000;
            14'h6571: o_data_a = 16'b1111000010001000;
            14'h6572: o_data_a = 16'b0000000000000000;
            14'h6573: o_data_a = 16'b1111110010101000;
            14'h6574: o_data_a = 16'b1111110000010000;
            14'h6575: o_data_a = 16'b0000000000000100;
            14'h6576: o_data_a = 16'b1110001100001000;
            14'h6577: o_data_a = 16'b0000000000000100;
            14'h6578: o_data_a = 16'b1111110000100000;
            14'h6579: o_data_a = 16'b1111110000010000;
            14'h657a: o_data_a = 16'b0000000000000000;
            14'h657b: o_data_a = 16'b1111110111101000;
            14'h657c: o_data_a = 16'b1110110010100000;
            14'h657d: o_data_a = 16'b1110001100001000;
            14'h657e: o_data_a = 16'b0000000000101101;
            14'h657f: o_data_a = 16'b1110110000010000;
            14'h6580: o_data_a = 16'b0000000000000000;
            14'h6581: o_data_a = 16'b1111110111101000;
            14'h6582: o_data_a = 16'b1110110010100000;
            14'h6583: o_data_a = 16'b1110001100001000;
            14'h6584: o_data_a = 16'b0110010110001000;
            14'h6585: o_data_a = 16'b1110110000010000;
            14'h6586: o_data_a = 16'b0000000000000110;
            14'h6587: o_data_a = 16'b1110101010000111;
            14'h6588: o_data_a = 16'b0000000000000000;
            14'h6589: o_data_a = 16'b1111110010101000;
            14'h658a: o_data_a = 16'b1111110000010000;
            14'h658b: o_data_a = 16'b0110010110001111;
            14'h658c: o_data_a = 16'b1110001100000101;
            14'h658d: o_data_a = 16'b0110010110101001;
            14'h658e: o_data_a = 16'b1110101010000111;
            14'h658f: o_data_a = 16'b0000000000000000;
            14'h6590: o_data_a = 16'b1111110111001000;
            14'h6591: o_data_a = 16'b1111110010100000;
            14'h6592: o_data_a = 16'b1110101010001000;
            14'h6593: o_data_a = 16'b0000000000000000;
            14'h6594: o_data_a = 16'b1111110010100000;
            14'h6595: o_data_a = 16'b1111110001001000;
            14'h6596: o_data_a = 16'b0000000000000000;
            14'h6597: o_data_a = 16'b1111110010101000;
            14'h6598: o_data_a = 16'b1111110000010000;
            14'h6599: o_data_a = 16'b0000000000000001;
            14'h659a: o_data_a = 16'b1111110111100000;
            14'h659b: o_data_a = 16'b1110110111100000;
            14'h659c: o_data_a = 16'b1110110111100000;
            14'h659d: o_data_a = 16'b1110110111100000;
            14'h659e: o_data_a = 16'b1110001100001000;
            14'h659f: o_data_a = 16'b0000000000000000;
            14'h65a0: o_data_a = 16'b1111110111001000;
            14'h65a1: o_data_a = 16'b1111110010100000;
            14'h65a2: o_data_a = 16'b1110111111001000;
            14'h65a3: o_data_a = 16'b0000000000000000;
            14'h65a4: o_data_a = 16'b1111110010101000;
            14'h65a5: o_data_a = 16'b1111110000010000;
            14'h65a6: o_data_a = 16'b0000000000000001;
            14'h65a7: o_data_a = 16'b1111110000100000;
            14'h65a8: o_data_a = 16'b1110001100001000;
            14'h65a9: o_data_a = 16'b0000000000000001;
            14'h65aa: o_data_a = 16'b1111110000100000;
            14'h65ab: o_data_a = 16'b1111110000010000;
            14'h65ac: o_data_a = 16'b0000000000000000;
            14'h65ad: o_data_a = 16'b1111110111101000;
            14'h65ae: o_data_a = 16'b1110110010100000;
            14'h65af: o_data_a = 16'b1110001100001000;
            14'h65b0: o_data_a = 16'b0000000000000011;
            14'h65b1: o_data_a = 16'b1111110111100000;
            14'h65b2: o_data_a = 16'b1110110111100000;
            14'h65b3: o_data_a = 16'b1111110000010000;
            14'h65b4: o_data_a = 16'b0000000000000000;
            14'h65b5: o_data_a = 16'b1111110111101000;
            14'h65b6: o_data_a = 16'b1110110010100000;
            14'h65b7: o_data_a = 16'b1110001100001000;
            14'h65b8: o_data_a = 16'b0110010110111100;
            14'h65b9: o_data_a = 16'b1110110000010000;
            14'h65ba: o_data_a = 16'b0000000000100110;
            14'h65bb: o_data_a = 16'b1110101010000111;
            14'h65bc: o_data_a = 16'b0000000000000001;
            14'h65bd: o_data_a = 16'b1111110000010000;
            14'h65be: o_data_a = 16'b0000000000000011;
            14'h65bf: o_data_a = 16'b1110000010100000;
            14'h65c0: o_data_a = 16'b1111110000010000;
            14'h65c1: o_data_a = 16'b0000000000000000;
            14'h65c2: o_data_a = 16'b1111110111101000;
            14'h65c3: o_data_a = 16'b1110110010100000;
            14'h65c4: o_data_a = 16'b1110001100001000;
            14'h65c5: o_data_a = 16'b0000000000000000;
            14'h65c6: o_data_a = 16'b1111110010101000;
            14'h65c7: o_data_a = 16'b1111110000010000;
            14'h65c8: o_data_a = 16'b1110110010100000;
            14'h65c9: o_data_a = 16'b1111000000001000;
            14'h65ca: o_data_a = 16'b0000000000000000;
            14'h65cb: o_data_a = 16'b1111110010100000;
            14'h65cc: o_data_a = 16'b1111110001001000;
            14'h65cd: o_data_a = 16'b0000000000000000;
            14'h65ce: o_data_a = 16'b1111110010101000;
            14'h65cf: o_data_a = 16'b1111110000010000;
            14'h65d0: o_data_a = 16'b0110011010001001;
            14'h65d1: o_data_a = 16'b1110001100000101;
            14'h65d2: o_data_a = 16'b0000000000000001;
            14'h65d3: o_data_a = 16'b1111110000100000;
            14'h65d4: o_data_a = 16'b1111110000010000;
            14'h65d5: o_data_a = 16'b0000000000000000;
            14'h65d6: o_data_a = 16'b1111110111101000;
            14'h65d7: o_data_a = 16'b1110110010100000;
            14'h65d8: o_data_a = 16'b1110001100001000;
            14'h65d9: o_data_a = 16'b0000000000000011;
            14'h65da: o_data_a = 16'b1111110111100000;
            14'h65db: o_data_a = 16'b1111110000010000;
            14'h65dc: o_data_a = 16'b0000000000000000;
            14'h65dd: o_data_a = 16'b1111110111101000;
            14'h65de: o_data_a = 16'b1110110010100000;
            14'h65df: o_data_a = 16'b1110001100001000;
            14'h65e0: o_data_a = 16'b0000000000000000;
            14'h65e1: o_data_a = 16'b1111110010101000;
            14'h65e2: o_data_a = 16'b1111110000010000;
            14'h65e3: o_data_a = 16'b1110110010100000;
            14'h65e4: o_data_a = 16'b1111000010001000;
            14'h65e5: o_data_a = 16'b0000000000000000;
            14'h65e6: o_data_a = 16'b1111110010101000;
            14'h65e7: o_data_a = 16'b1111110000010000;
            14'h65e8: o_data_a = 16'b0000000000000100;
            14'h65e9: o_data_a = 16'b1110001100001000;
            14'h65ea: o_data_a = 16'b0000000000000100;
            14'h65eb: o_data_a = 16'b1111110000100000;
            14'h65ec: o_data_a = 16'b1111110000010000;
            14'h65ed: o_data_a = 16'b0000000000000000;
            14'h65ee: o_data_a = 16'b1111110111101000;
            14'h65ef: o_data_a = 16'b1110110010100000;
            14'h65f0: o_data_a = 16'b1110001100001000;
            14'h65f1: o_data_a = 16'b0000000000110000;
            14'h65f2: o_data_a = 16'b1110110000010000;
            14'h65f3: o_data_a = 16'b0000000000000000;
            14'h65f4: o_data_a = 16'b1111110111101000;
            14'h65f5: o_data_a = 16'b1110110010100000;
            14'h65f6: o_data_a = 16'b1110001100001000;
            14'h65f7: o_data_a = 16'b0000000000000000;
            14'h65f8: o_data_a = 16'b1111110010101000;
            14'h65f9: o_data_a = 16'b1111110000010000;
            14'h65fa: o_data_a = 16'b1110110010100000;
            14'h65fb: o_data_a = 16'b1111000111001000;
            14'h65fc: o_data_a = 16'b0000000000000000;
            14'h65fd: o_data_a = 16'b1111110010101000;
            14'h65fe: o_data_a = 16'b1111110000010000;
            14'h65ff: o_data_a = 16'b0000000000000001;
            14'h6600: o_data_a = 16'b1111110111100000;
            14'h6601: o_data_a = 16'b1110110111100000;
            14'h6602: o_data_a = 16'b1110001100001000;
            14'h6603: o_data_a = 16'b0000000000000001;
            14'h6604: o_data_a = 16'b1111110111100000;
            14'h6605: o_data_a = 16'b1110110111100000;
            14'h6606: o_data_a = 16'b1111110000010000;
            14'h6607: o_data_a = 16'b0000000000000000;
            14'h6608: o_data_a = 16'b1111110111101000;
            14'h6609: o_data_a = 16'b1110110010100000;
            14'h660a: o_data_a = 16'b1110001100001000;
            14'h660b: o_data_a = 16'b0000000000000000;
            14'h660c: o_data_a = 16'b1111110111001000;
            14'h660d: o_data_a = 16'b1111110010100000;
            14'h660e: o_data_a = 16'b1110101010001000;
            14'h660f: o_data_a = 16'b0110011000010011;
            14'h6610: o_data_a = 16'b1110110000010000;
            14'h6611: o_data_a = 16'b0000000000100110;
            14'h6612: o_data_a = 16'b1110101010000111;
            14'h6613: o_data_a = 16'b0000000000000001;
            14'h6614: o_data_a = 16'b1111110111100000;
            14'h6615: o_data_a = 16'b1110110111100000;
            14'h6616: o_data_a = 16'b1111110000010000;
            14'h6617: o_data_a = 16'b0000000000000000;
            14'h6618: o_data_a = 16'b1111110111101000;
            14'h6619: o_data_a = 16'b1110110010100000;
            14'h661a: o_data_a = 16'b1110001100001000;
            14'h661b: o_data_a = 16'b0000000000001001;
            14'h661c: o_data_a = 16'b1110110000010000;
            14'h661d: o_data_a = 16'b0000000000000000;
            14'h661e: o_data_a = 16'b1111110111101000;
            14'h661f: o_data_a = 16'b1110110010100000;
            14'h6620: o_data_a = 16'b1110001100001000;
            14'h6621: o_data_a = 16'b0110011000100101;
            14'h6622: o_data_a = 16'b1110110000010000;
            14'h6623: o_data_a = 16'b0000000000010110;
            14'h6624: o_data_a = 16'b1110101010000111;
            14'h6625: o_data_a = 16'b0000000000000000;
            14'h6626: o_data_a = 16'b1111110010101000;
            14'h6627: o_data_a = 16'b1111110000010000;
            14'h6628: o_data_a = 16'b1110110010100000;
            14'h6629: o_data_a = 16'b1111010101001000;
            14'h662a: o_data_a = 16'b0000000000000000;
            14'h662b: o_data_a = 16'b1111110010100000;
            14'h662c: o_data_a = 16'b1111110001001000;
            14'h662d: o_data_a = 16'b0000000000000000;
            14'h662e: o_data_a = 16'b1111110010101000;
            14'h662f: o_data_a = 16'b1111110000010000;
            14'h6630: o_data_a = 16'b0000000000000001;
            14'h6631: o_data_a = 16'b1111110111100000;
            14'h6632: o_data_a = 16'b1110110111100000;
            14'h6633: o_data_a = 16'b1110110111100000;
            14'h6634: o_data_a = 16'b1110001100001000;
            14'h6635: o_data_a = 16'b0000000000000001;
            14'h6636: o_data_a = 16'b1111110000010000;
            14'h6637: o_data_a = 16'b0000000000000011;
            14'h6638: o_data_a = 16'b1110000010100000;
            14'h6639: o_data_a = 16'b1111110000010000;
            14'h663a: o_data_a = 16'b0000000000000000;
            14'h663b: o_data_a = 16'b1111110111101000;
            14'h663c: o_data_a = 16'b1110110010100000;
            14'h663d: o_data_a = 16'b1110001100001000;
            14'h663e: o_data_a = 16'b0000000000000000;
            14'h663f: o_data_a = 16'b1111110010101000;
            14'h6640: o_data_a = 16'b1111110000010000;
            14'h6641: o_data_a = 16'b0110011001000101;
            14'h6642: o_data_a = 16'b1110001100000101;
            14'h6643: o_data_a = 16'b0110011010000111;
            14'h6644: o_data_a = 16'b1110101010000111;
            14'h6645: o_data_a = 16'b0000000000000001;
            14'h6646: o_data_a = 16'b1111110111100000;
            14'h6647: o_data_a = 16'b1111110000010000;
            14'h6648: o_data_a = 16'b0000000000000000;
            14'h6649: o_data_a = 16'b1111110111101000;
            14'h664a: o_data_a = 16'b1110110010100000;
            14'h664b: o_data_a = 16'b1110001100001000;
            14'h664c: o_data_a = 16'b0000000000001010;
            14'h664d: o_data_a = 16'b1110110000010000;
            14'h664e: o_data_a = 16'b0000000000000000;
            14'h664f: o_data_a = 16'b1111110111101000;
            14'h6650: o_data_a = 16'b1110110010100000;
            14'h6651: o_data_a = 16'b1110001100001000;
            14'h6652: o_data_a = 16'b0000000000000010;
            14'h6653: o_data_a = 16'b1110110000010000;
            14'h6654: o_data_a = 16'b0000000000001101;
            14'h6655: o_data_a = 16'b1110001100001000;
            14'h6656: o_data_a = 16'b0001101010100110;
            14'h6657: o_data_a = 16'b1110110000010000;
            14'h6658: o_data_a = 16'b0000000000001110;
            14'h6659: o_data_a = 16'b1110001100001000;
            14'h665a: o_data_a = 16'b0110011001011110;
            14'h665b: o_data_a = 16'b1110110000010000;
            14'h665c: o_data_a = 16'b0000000001011111;
            14'h665d: o_data_a = 16'b1110101010000111;
            14'h665e: o_data_a = 16'b0000000000000001;
            14'h665f: o_data_a = 16'b1111110111100000;
            14'h6660: o_data_a = 16'b1110110111100000;
            14'h6661: o_data_a = 16'b1111110000010000;
            14'h6662: o_data_a = 16'b0000000000000000;
            14'h6663: o_data_a = 16'b1111110111101000;
            14'h6664: o_data_a = 16'b1110110010100000;
            14'h6665: o_data_a = 16'b1110001100001000;
            14'h6666: o_data_a = 16'b0000000000000000;
            14'h6667: o_data_a = 16'b1111110010101000;
            14'h6668: o_data_a = 16'b1111110000010000;
            14'h6669: o_data_a = 16'b1110110010100000;
            14'h666a: o_data_a = 16'b1111000010001000;
            14'h666b: o_data_a = 16'b0000000000000000;
            14'h666c: o_data_a = 16'b1111110010101000;
            14'h666d: o_data_a = 16'b1111110000010000;
            14'h666e: o_data_a = 16'b0000000000000001;
            14'h666f: o_data_a = 16'b1111110111100000;
            14'h6670: o_data_a = 16'b1110001100001000;
            14'h6671: o_data_a = 16'b0000000000000001;
            14'h6672: o_data_a = 16'b1111110000100000;
            14'h6673: o_data_a = 16'b1111110000010000;
            14'h6674: o_data_a = 16'b0000000000000000;
            14'h6675: o_data_a = 16'b1111110111101000;
            14'h6676: o_data_a = 16'b1110110010100000;
            14'h6677: o_data_a = 16'b1110001100001000;
            14'h6678: o_data_a = 16'b0000000000000000;
            14'h6679: o_data_a = 16'b1111110111001000;
            14'h667a: o_data_a = 16'b1111110010100000;
            14'h667b: o_data_a = 16'b1110111111001000;
            14'h667c: o_data_a = 16'b0000000000000000;
            14'h667d: o_data_a = 16'b1111110010101000;
            14'h667e: o_data_a = 16'b1111110000010000;
            14'h667f: o_data_a = 16'b1110110010100000;
            14'h6680: o_data_a = 16'b1111000010001000;
            14'h6681: o_data_a = 16'b0000000000000000;
            14'h6682: o_data_a = 16'b1111110010101000;
            14'h6683: o_data_a = 16'b1111110000010000;
            14'h6684: o_data_a = 16'b0000000000000001;
            14'h6685: o_data_a = 16'b1111110000100000;
            14'h6686: o_data_a = 16'b1110001100001000;
            14'h6687: o_data_a = 16'b0110010110101001;
            14'h6688: o_data_a = 16'b1110101010000111;
            14'h6689: o_data_a = 16'b0000000000000001;
            14'h668a: o_data_a = 16'b1111110000010000;
            14'h668b: o_data_a = 16'b0000000000000100;
            14'h668c: o_data_a = 16'b1110000010100000;
            14'h668d: o_data_a = 16'b1111110000010000;
            14'h668e: o_data_a = 16'b0000000000000000;
            14'h668f: o_data_a = 16'b1111110111101000;
            14'h6690: o_data_a = 16'b1110110010100000;
            14'h6691: o_data_a = 16'b1110001100001000;
            14'h6692: o_data_a = 16'b0000000000000000;
            14'h6693: o_data_a = 16'b1111110010101000;
            14'h6694: o_data_a = 16'b1111110000010000;
            14'h6695: o_data_a = 16'b0110011010011001;
            14'h6696: o_data_a = 16'b1110001100000101;
            14'h6697: o_data_a = 16'b0110011010101010;
            14'h6698: o_data_a = 16'b1110101010000111;
            14'h6699: o_data_a = 16'b0000000000000001;
            14'h669a: o_data_a = 16'b1111110111100000;
            14'h669b: o_data_a = 16'b1111110000010000;
            14'h669c: o_data_a = 16'b0000000000000000;
            14'h669d: o_data_a = 16'b1111110111101000;
            14'h669e: o_data_a = 16'b1110110010100000;
            14'h669f: o_data_a = 16'b1110001100001000;
            14'h66a0: o_data_a = 16'b0000000000000000;
            14'h66a1: o_data_a = 16'b1111110010100000;
            14'h66a2: o_data_a = 16'b1111110001010000;
            14'h66a3: o_data_a = 16'b1110011111001000;
            14'h66a4: o_data_a = 16'b0000000000000000;
            14'h66a5: o_data_a = 16'b1111110010101000;
            14'h66a6: o_data_a = 16'b1111110000010000;
            14'h66a7: o_data_a = 16'b0000000000000001;
            14'h66a8: o_data_a = 16'b1111110111100000;
            14'h66a9: o_data_a = 16'b1110001100001000;
            14'h66aa: o_data_a = 16'b0000000000000001;
            14'h66ab: o_data_a = 16'b1111110111100000;
            14'h66ac: o_data_a = 16'b1111110000010000;
            14'h66ad: o_data_a = 16'b0000000000000000;
            14'h66ae: o_data_a = 16'b1111110111101000;
            14'h66af: o_data_a = 16'b1110110010100000;
            14'h66b0: o_data_a = 16'b1110001100001000;
            14'h66b1: o_data_a = 16'b0000000000110110;
            14'h66b2: o_data_a = 16'b1110101010000111;
            14'h66b3: o_data_a = 16'b0000000000000100;
            14'h66b4: o_data_a = 16'b1110110000010000;
            14'h66b5: o_data_a = 16'b1110001110010000;
            14'h66b6: o_data_a = 16'b0000000000000000;
            14'h66b7: o_data_a = 16'b1111110111101000;
            14'h66b8: o_data_a = 16'b1110110010100000;
            14'h66b9: o_data_a = 16'b1110101010001000;
            14'h66ba: o_data_a = 16'b0110011010110101;
            14'h66bb: o_data_a = 16'b1110001100000001;
            14'h66bc: o_data_a = 16'b0000000000000010;
            14'h66bd: o_data_a = 16'b1111110000100000;
            14'h66be: o_data_a = 16'b1111110000010000;
            14'h66bf: o_data_a = 16'b0000000000000000;
            14'h66c0: o_data_a = 16'b1111110111101000;
            14'h66c1: o_data_a = 16'b1110110010100000;
            14'h66c2: o_data_a = 16'b1110001100001000;
            14'h66c3: o_data_a = 16'b0000000000000000;
            14'h66c4: o_data_a = 16'b1111110010101000;
            14'h66c5: o_data_a = 16'b1111110000010000;
            14'h66c6: o_data_a = 16'b0000000000000011;
            14'h66c7: o_data_a = 16'b1110001100001000;
            14'h66c8: o_data_a = 16'b0000000000000011;
            14'h66c9: o_data_a = 16'b1111110000100000;
            14'h66ca: o_data_a = 16'b1111110000010000;
            14'h66cb: o_data_a = 16'b0000000000000000;
            14'h66cc: o_data_a = 16'b1111110111101000;
            14'h66cd: o_data_a = 16'b1110110010100000;
            14'h66ce: o_data_a = 16'b1110001100001000;
            14'h66cf: o_data_a = 16'b0000000000000000;
            14'h66d0: o_data_a = 16'b1111110111001000;
            14'h66d1: o_data_a = 16'b1111110010100000;
            14'h66d2: o_data_a = 16'b1110101010001000;
            14'h66d3: o_data_a = 16'b0110011011010111;
            14'h66d4: o_data_a = 16'b1110110000010000;
            14'h66d5: o_data_a = 16'b0000000000000110;
            14'h66d6: o_data_a = 16'b1110101010000111;
            14'h66d7: o_data_a = 16'b0000000000000000;
            14'h66d8: o_data_a = 16'b1111110010101000;
            14'h66d9: o_data_a = 16'b1111110000010000;
            14'h66da: o_data_a = 16'b0110011011011110;
            14'h66db: o_data_a = 16'b1110001100000101;
            14'h66dc: o_data_a = 16'b0110011011110101;
            14'h66dd: o_data_a = 16'b1110101010000111;
            14'h66de: o_data_a = 16'b0000000000010011;
            14'h66df: o_data_a = 16'b1110110000010000;
            14'h66e0: o_data_a = 16'b0000000000000000;
            14'h66e1: o_data_a = 16'b1111110111101000;
            14'h66e2: o_data_a = 16'b1110110010100000;
            14'h66e3: o_data_a = 16'b1110001100001000;
            14'h66e4: o_data_a = 16'b0000000000000001;
            14'h66e5: o_data_a = 16'b1110110000010000;
            14'h66e6: o_data_a = 16'b0000000000001101;
            14'h66e7: o_data_a = 16'b1110001100001000;
            14'h66e8: o_data_a = 16'b0110101011011001;
            14'h66e9: o_data_a = 16'b1110110000010000;
            14'h66ea: o_data_a = 16'b0000000000001110;
            14'h66eb: o_data_a = 16'b1110001100001000;
            14'h66ec: o_data_a = 16'b0110011011110000;
            14'h66ed: o_data_a = 16'b1110110000010000;
            14'h66ee: o_data_a = 16'b0000000001011111;
            14'h66ef: o_data_a = 16'b1110101010000111;
            14'h66f0: o_data_a = 16'b0000000000000000;
            14'h66f1: o_data_a = 16'b1111110010101000;
            14'h66f2: o_data_a = 16'b1111110000010000;
            14'h66f3: o_data_a = 16'b0000000000000101;
            14'h66f4: o_data_a = 16'b1110001100001000;
            14'h66f5: o_data_a = 16'b0000000000000110;
            14'h66f6: o_data_a = 16'b1110110000010000;
            14'h66f7: o_data_a = 16'b0000000000000000;
            14'h66f8: o_data_a = 16'b1111110111101000;
            14'h66f9: o_data_a = 16'b1110110010100000;
            14'h66fa: o_data_a = 16'b1110001100001000;
            14'h66fb: o_data_a = 16'b0000000000000001;
            14'h66fc: o_data_a = 16'b1110110000010000;
            14'h66fd: o_data_a = 16'b0000000000001101;
            14'h66fe: o_data_a = 16'b1110001100001000;
            14'h66ff: o_data_a = 16'b0001011010110000;
            14'h6700: o_data_a = 16'b1110110000010000;
            14'h6701: o_data_a = 16'b0000000000001110;
            14'h6702: o_data_a = 16'b1110001100001000;
            14'h6703: o_data_a = 16'b0110011100000111;
            14'h6704: o_data_a = 16'b1110110000010000;
            14'h6705: o_data_a = 16'b0000000001011111;
            14'h6706: o_data_a = 16'b1110101010000111;
            14'h6707: o_data_a = 16'b0000000000000000;
            14'h6708: o_data_a = 16'b1111110010101000;
            14'h6709: o_data_a = 16'b1111110000010000;
            14'h670a: o_data_a = 16'b0000000000000001;
            14'h670b: o_data_a = 16'b1111110111100000;
            14'h670c: o_data_a = 16'b1110110111100000;
            14'h670d: o_data_a = 16'b1110001100001000;
            14'h670e: o_data_a = 16'b0000000000000010;
            14'h670f: o_data_a = 16'b1111110111100000;
            14'h6710: o_data_a = 16'b1111110000010000;
            14'h6711: o_data_a = 16'b0000000000000000;
            14'h6712: o_data_a = 16'b1111110111101000;
            14'h6713: o_data_a = 16'b1110110010100000;
            14'h6714: o_data_a = 16'b1110001100001000;
            14'h6715: o_data_a = 16'b0000000000000000;
            14'h6716: o_data_a = 16'b1111110111001000;
            14'h6717: o_data_a = 16'b1111110010100000;
            14'h6718: o_data_a = 16'b1110101010001000;
            14'h6719: o_data_a = 16'b0110011100011101;
            14'h671a: o_data_a = 16'b1110110000010000;
            14'h671b: o_data_a = 16'b0000000000100110;
            14'h671c: o_data_a = 16'b1110101010000111;
            14'h671d: o_data_a = 16'b0000000000000000;
            14'h671e: o_data_a = 16'b1111110010101000;
            14'h671f: o_data_a = 16'b1111110000010000;
            14'h6720: o_data_a = 16'b0110011100100100;
            14'h6721: o_data_a = 16'b1110001100000101;
            14'h6722: o_data_a = 16'b0110011101000100;
            14'h6723: o_data_a = 16'b1110101010000111;
            14'h6724: o_data_a = 16'b0000000000000000;
            14'h6725: o_data_a = 16'b1111110111001000;
            14'h6726: o_data_a = 16'b1111110010100000;
            14'h6727: o_data_a = 16'b1110101010001000;
            14'h6728: o_data_a = 16'b0000000000000000;
            14'h6729: o_data_a = 16'b1111110010100000;
            14'h672a: o_data_a = 16'b1111110001001000;
            14'h672b: o_data_a = 16'b0000000000000000;
            14'h672c: o_data_a = 16'b1111110010101000;
            14'h672d: o_data_a = 16'b1111110000010000;
            14'h672e: o_data_a = 16'b0000000000000001;
            14'h672f: o_data_a = 16'b1111110111100000;
            14'h6730: o_data_a = 16'b1110110111100000;
            14'h6731: o_data_a = 16'b1110110111100000;
            14'h6732: o_data_a = 16'b1110001100001000;
            14'h6733: o_data_a = 16'b0000000000000010;
            14'h6734: o_data_a = 16'b1111110111100000;
            14'h6735: o_data_a = 16'b1111110000010000;
            14'h6736: o_data_a = 16'b0000000000000000;
            14'h6737: o_data_a = 16'b1111110111101000;
            14'h6738: o_data_a = 16'b1110110010100000;
            14'h6739: o_data_a = 16'b1110001100001000;
            14'h673a: o_data_a = 16'b0000000000000000;
            14'h673b: o_data_a = 16'b1111110010100000;
            14'h673c: o_data_a = 16'b1111110001010000;
            14'h673d: o_data_a = 16'b1110011111001000;
            14'h673e: o_data_a = 16'b0000000000000000;
            14'h673f: o_data_a = 16'b1111110010101000;
            14'h6740: o_data_a = 16'b1111110000010000;
            14'h6741: o_data_a = 16'b0000000000000010;
            14'h6742: o_data_a = 16'b1111110111100000;
            14'h6743: o_data_a = 16'b1110001100001000;
            14'h6744: o_data_a = 16'b0000000000000010;
            14'h6745: o_data_a = 16'b1111110111100000;
            14'h6746: o_data_a = 16'b1111110000010000;
            14'h6747: o_data_a = 16'b0000000000000000;
            14'h6748: o_data_a = 16'b1111110111101000;
            14'h6749: o_data_a = 16'b1110110010100000;
            14'h674a: o_data_a = 16'b1110001100001000;
            14'h674b: o_data_a = 16'b0000000000000000;
            14'h674c: o_data_a = 16'b1111110010101000;
            14'h674d: o_data_a = 16'b1111110000010000;
            14'h674e: o_data_a = 16'b0000000000000001;
            14'h674f: o_data_a = 16'b1111110111100000;
            14'h6750: o_data_a = 16'b1110001100001000;
            14'h6751: o_data_a = 16'b0000000000000001;
            14'h6752: o_data_a = 16'b1111110111100000;
            14'h6753: o_data_a = 16'b1111110000010000;
            14'h6754: o_data_a = 16'b0000000000000000;
            14'h6755: o_data_a = 16'b1111110111101000;
            14'h6756: o_data_a = 16'b1110110010100000;
            14'h6757: o_data_a = 16'b1110001100001000;
            14'h6758: o_data_a = 16'b0000000000000000;
            14'h6759: o_data_a = 16'b1111110111001000;
            14'h675a: o_data_a = 16'b1111110010100000;
            14'h675b: o_data_a = 16'b1110101010001000;
            14'h675c: o_data_a = 16'b0110011101100000;
            14'h675d: o_data_a = 16'b1110110000010000;
            14'h675e: o_data_a = 16'b0000000000010110;
            14'h675f: o_data_a = 16'b1110101010000111;
            14'h6760: o_data_a = 16'b0000000000000000;
            14'h6761: o_data_a = 16'b1111110010100000;
            14'h6762: o_data_a = 16'b1111110001001000;
            14'h6763: o_data_a = 16'b0000000000000000;
            14'h6764: o_data_a = 16'b1111110010101000;
            14'h6765: o_data_a = 16'b1111110000010000;
            14'h6766: o_data_a = 16'b0110100000000110;
            14'h6767: o_data_a = 16'b1110001100000101;
            14'h6768: o_data_a = 16'b0000000000000010;
            14'h6769: o_data_a = 16'b1111110111100000;
            14'h676a: o_data_a = 16'b1111110000010000;
            14'h676b: o_data_a = 16'b0000000000000000;
            14'h676c: o_data_a = 16'b1111110111101000;
            14'h676d: o_data_a = 16'b1110110010100000;
            14'h676e: o_data_a = 16'b1110001100001000;
            14'h676f: o_data_a = 16'b0000000000001010;
            14'h6770: o_data_a = 16'b1110110000010000;
            14'h6771: o_data_a = 16'b0000000000000000;
            14'h6772: o_data_a = 16'b1111110111101000;
            14'h6773: o_data_a = 16'b1110110010100000;
            14'h6774: o_data_a = 16'b1110001100001000;
            14'h6775: o_data_a = 16'b0000000000000010;
            14'h6776: o_data_a = 16'b1110110000010000;
            14'h6777: o_data_a = 16'b0000000000001101;
            14'h6778: o_data_a = 16'b1110001100001000;
            14'h6779: o_data_a = 16'b0001110001110111;
            14'h677a: o_data_a = 16'b1110110000010000;
            14'h677b: o_data_a = 16'b0000000000001110;
            14'h677c: o_data_a = 16'b1110001100001000;
            14'h677d: o_data_a = 16'b0110011110000001;
            14'h677e: o_data_a = 16'b1110110000010000;
            14'h677f: o_data_a = 16'b0000000001011111;
            14'h6780: o_data_a = 16'b1110101010000111;
            14'h6781: o_data_a = 16'b0000000000000000;
            14'h6782: o_data_a = 16'b1111110010101000;
            14'h6783: o_data_a = 16'b1111110000010000;
            14'h6784: o_data_a = 16'b0000000000000001;
            14'h6785: o_data_a = 16'b1111110111100000;
            14'h6786: o_data_a = 16'b1110001100001000;
            14'h6787: o_data_a = 16'b0000000000000001;
            14'h6788: o_data_a = 16'b1111110000100000;
            14'h6789: o_data_a = 16'b1111110000010000;
            14'h678a: o_data_a = 16'b0000000000000000;
            14'h678b: o_data_a = 16'b1111110111101000;
            14'h678c: o_data_a = 16'b1110110010100000;
            14'h678d: o_data_a = 16'b1110001100001000;
            14'h678e: o_data_a = 16'b0000000000000001;
            14'h678f: o_data_a = 16'b1111110111100000;
            14'h6790: o_data_a = 16'b1110110111100000;
            14'h6791: o_data_a = 16'b1111110000010000;
            14'h6792: o_data_a = 16'b0000000000000000;
            14'h6793: o_data_a = 16'b1111110111101000;
            14'h6794: o_data_a = 16'b1110110010100000;
            14'h6795: o_data_a = 16'b1110001100001000;
            14'h6796: o_data_a = 16'b0000000000000000;
            14'h6797: o_data_a = 16'b1111110010101000;
            14'h6798: o_data_a = 16'b1111110000010000;
            14'h6799: o_data_a = 16'b1110110010100000;
            14'h679a: o_data_a = 16'b1111000010001000;
            14'h679b: o_data_a = 16'b0000000000110000;
            14'h679c: o_data_a = 16'b1110110000010000;
            14'h679d: o_data_a = 16'b0000000000000000;
            14'h679e: o_data_a = 16'b1111110111101000;
            14'h679f: o_data_a = 16'b1110110010100000;
            14'h67a0: o_data_a = 16'b1110001100001000;
            14'h67a1: o_data_a = 16'b0000000000000010;
            14'h67a2: o_data_a = 16'b1111110111100000;
            14'h67a3: o_data_a = 16'b1111110000010000;
            14'h67a4: o_data_a = 16'b0000000000000000;
            14'h67a5: o_data_a = 16'b1111110111101000;
            14'h67a6: o_data_a = 16'b1110110010100000;
            14'h67a7: o_data_a = 16'b1110001100001000;
            14'h67a8: o_data_a = 16'b0000000000000001;
            14'h67a9: o_data_a = 16'b1111110111100000;
            14'h67aa: o_data_a = 16'b1111110000010000;
            14'h67ab: o_data_a = 16'b0000000000000000;
            14'h67ac: o_data_a = 16'b1111110111101000;
            14'h67ad: o_data_a = 16'b1110110010100000;
            14'h67ae: o_data_a = 16'b1110001100001000;
            14'h67af: o_data_a = 16'b0000000000001010;
            14'h67b0: o_data_a = 16'b1110110000010000;
            14'h67b1: o_data_a = 16'b0000000000000000;
            14'h67b2: o_data_a = 16'b1111110111101000;
            14'h67b3: o_data_a = 16'b1110110010100000;
            14'h67b4: o_data_a = 16'b1110001100001000;
            14'h67b5: o_data_a = 16'b0000000000000010;
            14'h67b6: o_data_a = 16'b1110110000010000;
            14'h67b7: o_data_a = 16'b0000000000001101;
            14'h67b8: o_data_a = 16'b1110001100001000;
            14'h67b9: o_data_a = 16'b0001101010100110;
            14'h67ba: o_data_a = 16'b1110110000010000;
            14'h67bb: o_data_a = 16'b0000000000001110;
            14'h67bc: o_data_a = 16'b1110001100001000;
            14'h67bd: o_data_a = 16'b0110011111000001;
            14'h67be: o_data_a = 16'b1110110000010000;
            14'h67bf: o_data_a = 16'b0000000001011111;
            14'h67c0: o_data_a = 16'b1110101010000111;
            14'h67c1: o_data_a = 16'b0000000000000000;
            14'h67c2: o_data_a = 16'b1111110010101000;
            14'h67c3: o_data_a = 16'b1111110000010000;
            14'h67c4: o_data_a = 16'b1110110010100000;
            14'h67c5: o_data_a = 16'b1111000111001000;
            14'h67c6: o_data_a = 16'b0000000000000000;
            14'h67c7: o_data_a = 16'b1111110010101000;
            14'h67c8: o_data_a = 16'b1111110000010000;
            14'h67c9: o_data_a = 16'b1110110010100000;
            14'h67ca: o_data_a = 16'b1111000010001000;
            14'h67cb: o_data_a = 16'b0000000000000000;
            14'h67cc: o_data_a = 16'b1111110010101000;
            14'h67cd: o_data_a = 16'b1111110000010000;
            14'h67ce: o_data_a = 16'b0000000000000101;
            14'h67cf: o_data_a = 16'b1110001100001000;
            14'h67d0: o_data_a = 16'b0000000000000000;
            14'h67d1: o_data_a = 16'b1111110010101000;
            14'h67d2: o_data_a = 16'b1111110000010000;
            14'h67d3: o_data_a = 16'b0000000000000100;
            14'h67d4: o_data_a = 16'b1110001100001000;
            14'h67d5: o_data_a = 16'b0000000000000101;
            14'h67d6: o_data_a = 16'b1111110000010000;
            14'h67d7: o_data_a = 16'b0000000000000000;
            14'h67d8: o_data_a = 16'b1111110111101000;
            14'h67d9: o_data_a = 16'b1110110010100000;
            14'h67da: o_data_a = 16'b1110001100001000;
            14'h67db: o_data_a = 16'b0000000000000000;
            14'h67dc: o_data_a = 16'b1111110010101000;
            14'h67dd: o_data_a = 16'b1111110000010000;
            14'h67de: o_data_a = 16'b0000000000000100;
            14'h67df: o_data_a = 16'b1111110000100000;
            14'h67e0: o_data_a = 16'b1110001100001000;
            14'h67e1: o_data_a = 16'b0000000000000001;
            14'h67e2: o_data_a = 16'b1111110000100000;
            14'h67e3: o_data_a = 16'b1111110000010000;
            14'h67e4: o_data_a = 16'b0000000000000000;
            14'h67e5: o_data_a = 16'b1111110111101000;
            14'h67e6: o_data_a = 16'b1110110010100000;
            14'h67e7: o_data_a = 16'b1110001100001000;
            14'h67e8: o_data_a = 16'b0000000000000000;
            14'h67e9: o_data_a = 16'b1111110111001000;
            14'h67ea: o_data_a = 16'b1111110010100000;
            14'h67eb: o_data_a = 16'b1110111111001000;
            14'h67ec: o_data_a = 16'b0000000000000000;
            14'h67ed: o_data_a = 16'b1111110010101000;
            14'h67ee: o_data_a = 16'b1111110000010000;
            14'h67ef: o_data_a = 16'b1110110010100000;
            14'h67f0: o_data_a = 16'b1111000010001000;
            14'h67f1: o_data_a = 16'b0000000000000000;
            14'h67f2: o_data_a = 16'b1111110010101000;
            14'h67f3: o_data_a = 16'b1111110000010000;
            14'h67f4: o_data_a = 16'b0000000000000001;
            14'h67f5: o_data_a = 16'b1111110000100000;
            14'h67f6: o_data_a = 16'b1110001100001000;
            14'h67f7: o_data_a = 16'b0000000000000001;
            14'h67f8: o_data_a = 16'b1111110111100000;
            14'h67f9: o_data_a = 16'b1111110000010000;
            14'h67fa: o_data_a = 16'b0000000000000000;
            14'h67fb: o_data_a = 16'b1111110111101000;
            14'h67fc: o_data_a = 16'b1110110010100000;
            14'h67fd: o_data_a = 16'b1110001100001000;
            14'h67fe: o_data_a = 16'b0000000000000000;
            14'h67ff: o_data_a = 16'b1111110010101000;
            14'h6800: o_data_a = 16'b1111110000010000;
            14'h6801: o_data_a = 16'b0000000000000010;
            14'h6802: o_data_a = 16'b1111110111100000;
            14'h6803: o_data_a = 16'b1110001100001000;
            14'h6804: o_data_a = 16'b0110011101010001;
            14'h6805: o_data_a = 16'b1110101010000111;
            14'h6806: o_data_a = 16'b0000000000000001;
            14'h6807: o_data_a = 16'b1111110000010000;
            14'h6808: o_data_a = 16'b0000000000000011;
            14'h6809: o_data_a = 16'b1110000010100000;
            14'h680a: o_data_a = 16'b1111110000010000;
            14'h680b: o_data_a = 16'b0000000000000000;
            14'h680c: o_data_a = 16'b1111110111101000;
            14'h680d: o_data_a = 16'b1110110010100000;
            14'h680e: o_data_a = 16'b1110001100001000;
            14'h680f: o_data_a = 16'b0000000000000000;
            14'h6810: o_data_a = 16'b1111110010101000;
            14'h6811: o_data_a = 16'b1111110000010000;
            14'h6812: o_data_a = 16'b0110100000010110;
            14'h6813: o_data_a = 16'b1110001100000101;
            14'h6814: o_data_a = 16'b0110100001011100;
            14'h6815: o_data_a = 16'b1110101010000111;
            14'h6816: o_data_a = 16'b0000000000000001;
            14'h6817: o_data_a = 16'b1111110000100000;
            14'h6818: o_data_a = 16'b1111110000010000;
            14'h6819: o_data_a = 16'b0000000000000000;
            14'h681a: o_data_a = 16'b1111110111101000;
            14'h681b: o_data_a = 16'b1110110010100000;
            14'h681c: o_data_a = 16'b1110001100001000;
            14'h681d: o_data_a = 16'b0000000000000001;
            14'h681e: o_data_a = 16'b1111110111100000;
            14'h681f: o_data_a = 16'b1110110111100000;
            14'h6820: o_data_a = 16'b1111110000010000;
            14'h6821: o_data_a = 16'b0000000000000000;
            14'h6822: o_data_a = 16'b1111110111101000;
            14'h6823: o_data_a = 16'b1110110010100000;
            14'h6824: o_data_a = 16'b1110001100001000;
            14'h6825: o_data_a = 16'b0000000000000000;
            14'h6826: o_data_a = 16'b1111110010101000;
            14'h6827: o_data_a = 16'b1111110000010000;
            14'h6828: o_data_a = 16'b1110110010100000;
            14'h6829: o_data_a = 16'b1111000010001000;
            14'h682a: o_data_a = 16'b0000000000101101;
            14'h682b: o_data_a = 16'b1110110000010000;
            14'h682c: o_data_a = 16'b0000000000000000;
            14'h682d: o_data_a = 16'b1111110111101000;
            14'h682e: o_data_a = 16'b1110110010100000;
            14'h682f: o_data_a = 16'b1110001100001000;
            14'h6830: o_data_a = 16'b0000000000000000;
            14'h6831: o_data_a = 16'b1111110010101000;
            14'h6832: o_data_a = 16'b1111110000010000;
            14'h6833: o_data_a = 16'b0000000000000101;
            14'h6834: o_data_a = 16'b1110001100001000;
            14'h6835: o_data_a = 16'b0000000000000000;
            14'h6836: o_data_a = 16'b1111110010101000;
            14'h6837: o_data_a = 16'b1111110000010000;
            14'h6838: o_data_a = 16'b0000000000000100;
            14'h6839: o_data_a = 16'b1110001100001000;
            14'h683a: o_data_a = 16'b0000000000000101;
            14'h683b: o_data_a = 16'b1111110000010000;
            14'h683c: o_data_a = 16'b0000000000000000;
            14'h683d: o_data_a = 16'b1111110111101000;
            14'h683e: o_data_a = 16'b1110110010100000;
            14'h683f: o_data_a = 16'b1110001100001000;
            14'h6840: o_data_a = 16'b0000000000000000;
            14'h6841: o_data_a = 16'b1111110010101000;
            14'h6842: o_data_a = 16'b1111110000010000;
            14'h6843: o_data_a = 16'b0000000000000100;
            14'h6844: o_data_a = 16'b1111110000100000;
            14'h6845: o_data_a = 16'b1110001100001000;
            14'h6846: o_data_a = 16'b0000000000000001;
            14'h6847: o_data_a = 16'b1111110000100000;
            14'h6848: o_data_a = 16'b1111110000010000;
            14'h6849: o_data_a = 16'b0000000000000000;
            14'h684a: o_data_a = 16'b1111110111101000;
            14'h684b: o_data_a = 16'b1110110010100000;
            14'h684c: o_data_a = 16'b1110001100001000;
            14'h684d: o_data_a = 16'b0000000000000000;
            14'h684e: o_data_a = 16'b1111110111001000;
            14'h684f: o_data_a = 16'b1111110010100000;
            14'h6850: o_data_a = 16'b1110111111001000;
            14'h6851: o_data_a = 16'b0000000000000000;
            14'h6852: o_data_a = 16'b1111110010101000;
            14'h6853: o_data_a = 16'b1111110000010000;
            14'h6854: o_data_a = 16'b1110110010100000;
            14'h6855: o_data_a = 16'b1111000010001000;
            14'h6856: o_data_a = 16'b0000000000000000;
            14'h6857: o_data_a = 16'b1111110010101000;
            14'h6858: o_data_a = 16'b1111110000010000;
            14'h6859: o_data_a = 16'b0000000000000001;
            14'h685a: o_data_a = 16'b1111110000100000;
            14'h685b: o_data_a = 16'b1110001100001000;
            14'h685c: o_data_a = 16'b0000000000000011;
            14'h685d: o_data_a = 16'b1111110000100000;
            14'h685e: o_data_a = 16'b1111110000010000;
            14'h685f: o_data_a = 16'b0000000000000000;
            14'h6860: o_data_a = 16'b1111110111101000;
            14'h6861: o_data_a = 16'b1110110010100000;
            14'h6862: o_data_a = 16'b1110001100001000;
            14'h6863: o_data_a = 16'b0000000000000001;
            14'h6864: o_data_a = 16'b1111110000100000;
            14'h6865: o_data_a = 16'b1111110000010000;
            14'h6866: o_data_a = 16'b0000000000000000;
            14'h6867: o_data_a = 16'b1111110111101000;
            14'h6868: o_data_a = 16'b1110110010100000;
            14'h6869: o_data_a = 16'b1110001100001000;
            14'h686a: o_data_a = 16'b0110100001101110;
            14'h686b: o_data_a = 16'b1110110000010000;
            14'h686c: o_data_a = 16'b0000000000100110;
            14'h686d: o_data_a = 16'b1110101010000111;
            14'h686e: o_data_a = 16'b0000000000000000;
            14'h686f: o_data_a = 16'b1111110010101000;
            14'h6870: o_data_a = 16'b1111110000010000;
            14'h6871: o_data_a = 16'b0110100001110101;
            14'h6872: o_data_a = 16'b1110001100000101;
            14'h6873: o_data_a = 16'b0110100010001100;
            14'h6874: o_data_a = 16'b1110101010000111;
            14'h6875: o_data_a = 16'b0000000000010011;
            14'h6876: o_data_a = 16'b1110110000010000;
            14'h6877: o_data_a = 16'b0000000000000000;
            14'h6878: o_data_a = 16'b1111110111101000;
            14'h6879: o_data_a = 16'b1110110010100000;
            14'h687a: o_data_a = 16'b1110001100001000;
            14'h687b: o_data_a = 16'b0000000000000001;
            14'h687c: o_data_a = 16'b1110110000010000;
            14'h687d: o_data_a = 16'b0000000000001101;
            14'h687e: o_data_a = 16'b1110001100001000;
            14'h687f: o_data_a = 16'b0110101011011001;
            14'h6880: o_data_a = 16'b1110110000010000;
            14'h6881: o_data_a = 16'b0000000000001110;
            14'h6882: o_data_a = 16'b1110001100001000;
            14'h6883: o_data_a = 16'b0110100010000111;
            14'h6884: o_data_a = 16'b1110110000010000;
            14'h6885: o_data_a = 16'b0000000001011111;
            14'h6886: o_data_a = 16'b1110101010000111;
            14'h6887: o_data_a = 16'b0000000000000000;
            14'h6888: o_data_a = 16'b1111110010101000;
            14'h6889: o_data_a = 16'b1111110000010000;
            14'h688a: o_data_a = 16'b0000000000000101;
            14'h688b: o_data_a = 16'b1110001100001000;
            14'h688c: o_data_a = 16'b0000000000000001;
            14'h688d: o_data_a = 16'b1111110000100000;
            14'h688e: o_data_a = 16'b1111110000010000;
            14'h688f: o_data_a = 16'b0000000000000000;
            14'h6890: o_data_a = 16'b1111110111101000;
            14'h6891: o_data_a = 16'b1110110010100000;
            14'h6892: o_data_a = 16'b1110001100001000;
            14'h6893: o_data_a = 16'b0000000000000000;
            14'h6894: o_data_a = 16'b1111110111001000;
            14'h6895: o_data_a = 16'b1111110010100000;
            14'h6896: o_data_a = 16'b1110101010001000;
            14'h6897: o_data_a = 16'b0110100010011011;
            14'h6898: o_data_a = 16'b1110110000010000;
            14'h6899: o_data_a = 16'b0000000000000110;
            14'h689a: o_data_a = 16'b1110101010000111;
            14'h689b: o_data_a = 16'b0000000000000000;
            14'h689c: o_data_a = 16'b1111110010101000;
            14'h689d: o_data_a = 16'b1111110000010000;
            14'h689e: o_data_a = 16'b0110100010100010;
            14'h689f: o_data_a = 16'b1110001100000101;
            14'h68a0: o_data_a = 16'b0110100011011011;
            14'h68a1: o_data_a = 16'b1110101010000111;
            14'h68a2: o_data_a = 16'b0000000000000000;
            14'h68a3: o_data_a = 16'b1111110111001000;
            14'h68a4: o_data_a = 16'b1111110010100000;
            14'h68a5: o_data_a = 16'b1110101010001000;
            14'h68a6: o_data_a = 16'b0000000000000011;
            14'h68a7: o_data_a = 16'b1111110111100000;
            14'h68a8: o_data_a = 16'b1111110000010000;
            14'h68a9: o_data_a = 16'b0000000000000000;
            14'h68aa: o_data_a = 16'b1111110111101000;
            14'h68ab: o_data_a = 16'b1110110010100000;
            14'h68ac: o_data_a = 16'b1110001100001000;
            14'h68ad: o_data_a = 16'b0000000000000000;
            14'h68ae: o_data_a = 16'b1111110010101000;
            14'h68af: o_data_a = 16'b1111110000010000;
            14'h68b0: o_data_a = 16'b1110110010100000;
            14'h68b1: o_data_a = 16'b1111000010001000;
            14'h68b2: o_data_a = 16'b0000000000110000;
            14'h68b3: o_data_a = 16'b1110110000010000;
            14'h68b4: o_data_a = 16'b0000000000000000;
            14'h68b5: o_data_a = 16'b1111110111101000;
            14'h68b6: o_data_a = 16'b1110110010100000;
            14'h68b7: o_data_a = 16'b1110001100001000;
            14'h68b8: o_data_a = 16'b0000000000000000;
            14'h68b9: o_data_a = 16'b1111110010101000;
            14'h68ba: o_data_a = 16'b1111110000010000;
            14'h68bb: o_data_a = 16'b0000000000000101;
            14'h68bc: o_data_a = 16'b1110001100001000;
            14'h68bd: o_data_a = 16'b0000000000000000;
            14'h68be: o_data_a = 16'b1111110010101000;
            14'h68bf: o_data_a = 16'b1111110000010000;
            14'h68c0: o_data_a = 16'b0000000000000100;
            14'h68c1: o_data_a = 16'b1110001100001000;
            14'h68c2: o_data_a = 16'b0000000000000101;
            14'h68c3: o_data_a = 16'b1111110000010000;
            14'h68c4: o_data_a = 16'b0000000000000000;
            14'h68c5: o_data_a = 16'b1111110111101000;
            14'h68c6: o_data_a = 16'b1110110010100000;
            14'h68c7: o_data_a = 16'b1110001100001000;
            14'h68c8: o_data_a = 16'b0000000000000000;
            14'h68c9: o_data_a = 16'b1111110010101000;
            14'h68ca: o_data_a = 16'b1111110000010000;
            14'h68cb: o_data_a = 16'b0000000000000100;
            14'h68cc: o_data_a = 16'b1111110000100000;
            14'h68cd: o_data_a = 16'b1110001100001000;
            14'h68ce: o_data_a = 16'b0000000000000000;
            14'h68cf: o_data_a = 16'b1111110111001000;
            14'h68d0: o_data_a = 16'b1111110010100000;
            14'h68d1: o_data_a = 16'b1110111111001000;
            14'h68d2: o_data_a = 16'b0000000000000000;
            14'h68d3: o_data_a = 16'b1111110010101000;
            14'h68d4: o_data_a = 16'b1111110000010000;
            14'h68d5: o_data_a = 16'b0000000000000011;
            14'h68d6: o_data_a = 16'b1111110111100000;
            14'h68d7: o_data_a = 16'b1110110111100000;
            14'h68d8: o_data_a = 16'b1110001100001000;
            14'h68d9: o_data_a = 16'b0110100101111011;
            14'h68da: o_data_a = 16'b1110101010000111;
            14'h68db: o_data_a = 16'b0000000000000000;
            14'h68dc: o_data_a = 16'b1111110111001000;
            14'h68dd: o_data_a = 16'b1111110010100000;
            14'h68de: o_data_a = 16'b1110101010001000;
            14'h68df: o_data_a = 16'b0000000000000000;
            14'h68e0: o_data_a = 16'b1111110010101000;
            14'h68e1: o_data_a = 16'b1111110000010000;
            14'h68e2: o_data_a = 16'b0000000000000011;
            14'h68e3: o_data_a = 16'b1111110111100000;
            14'h68e4: o_data_a = 16'b1110110111100000;
            14'h68e5: o_data_a = 16'b1110001100001000;
            14'h68e6: o_data_a = 16'b0000000000000011;
            14'h68e7: o_data_a = 16'b1111110111100000;
            14'h68e8: o_data_a = 16'b1110110111100000;
            14'h68e9: o_data_a = 16'b1111110000010000;
            14'h68ea: o_data_a = 16'b0000000000000000;
            14'h68eb: o_data_a = 16'b1111110111101000;
            14'h68ec: o_data_a = 16'b1110110010100000;
            14'h68ed: o_data_a = 16'b1110001100001000;
            14'h68ee: o_data_a = 16'b0000000000000001;
            14'h68ef: o_data_a = 16'b1111110000100000;
            14'h68f0: o_data_a = 16'b1111110000010000;
            14'h68f1: o_data_a = 16'b0000000000000000;
            14'h68f2: o_data_a = 16'b1111110111101000;
            14'h68f3: o_data_a = 16'b1110110010100000;
            14'h68f4: o_data_a = 16'b1110001100001000;
            14'h68f5: o_data_a = 16'b0110100011111001;
            14'h68f6: o_data_a = 16'b1110110000010000;
            14'h68f7: o_data_a = 16'b0000000000100110;
            14'h68f8: o_data_a = 16'b1110101010000111;
            14'h68f9: o_data_a = 16'b0000000000000000;
            14'h68fa: o_data_a = 16'b1111110010100000;
            14'h68fb: o_data_a = 16'b1111110001001000;
            14'h68fc: o_data_a = 16'b0000000000000000;
            14'h68fd: o_data_a = 16'b1111110010101000;
            14'h68fe: o_data_a = 16'b1111110000010000;
            14'h68ff: o_data_a = 16'b0110100101111011;
            14'h6900: o_data_a = 16'b1110001100000101;
            14'h6901: o_data_a = 16'b0000000000000011;
            14'h6902: o_data_a = 16'b1111110111100000;
            14'h6903: o_data_a = 16'b1110110111100000;
            14'h6904: o_data_a = 16'b1111110000010000;
            14'h6905: o_data_a = 16'b0000000000000000;
            14'h6906: o_data_a = 16'b1111110111101000;
            14'h6907: o_data_a = 16'b1110110010100000;
            14'h6908: o_data_a = 16'b1110001100001000;
            14'h6909: o_data_a = 16'b0000000000000011;
            14'h690a: o_data_a = 16'b1111110111100000;
            14'h690b: o_data_a = 16'b1111110000010000;
            14'h690c: o_data_a = 16'b0000000000000000;
            14'h690d: o_data_a = 16'b1111110111101000;
            14'h690e: o_data_a = 16'b1110110010100000;
            14'h690f: o_data_a = 16'b1110001100001000;
            14'h6910: o_data_a = 16'b0000000000000000;
            14'h6911: o_data_a = 16'b1111110010101000;
            14'h6912: o_data_a = 16'b1111110000010000;
            14'h6913: o_data_a = 16'b1110110010100000;
            14'h6914: o_data_a = 16'b1111000010001000;
            14'h6915: o_data_a = 16'b0000000000000001;
            14'h6916: o_data_a = 16'b1111110000100000;
            14'h6917: o_data_a = 16'b1111110000010000;
            14'h6918: o_data_a = 16'b0000000000000000;
            14'h6919: o_data_a = 16'b1111110111101000;
            14'h691a: o_data_a = 16'b1110110010100000;
            14'h691b: o_data_a = 16'b1110001100001000;
            14'h691c: o_data_a = 16'b0000000000000011;
            14'h691d: o_data_a = 16'b1111110111100000;
            14'h691e: o_data_a = 16'b1110110111100000;
            14'h691f: o_data_a = 16'b1111110000010000;
            14'h6920: o_data_a = 16'b0000000000000000;
            14'h6921: o_data_a = 16'b1111110111101000;
            14'h6922: o_data_a = 16'b1110110010100000;
            14'h6923: o_data_a = 16'b1110001100001000;
            14'h6924: o_data_a = 16'b0000000000000000;
            14'h6925: o_data_a = 16'b1111110111001000;
            14'h6926: o_data_a = 16'b1111110010100000;
            14'h6927: o_data_a = 16'b1110111111001000;
            14'h6928: o_data_a = 16'b0000000000000000;
            14'h6929: o_data_a = 16'b1111110010101000;
            14'h692a: o_data_a = 16'b1111110000010000;
            14'h692b: o_data_a = 16'b1110110010100000;
            14'h692c: o_data_a = 16'b1111000010001000;
            14'h692d: o_data_a = 16'b0000000000000000;
            14'h692e: o_data_a = 16'b1111110010101000;
            14'h692f: o_data_a = 16'b1111110000010000;
            14'h6930: o_data_a = 16'b1110110010100000;
            14'h6931: o_data_a = 16'b1111000111001000;
            14'h6932: o_data_a = 16'b0000000000000001;
            14'h6933: o_data_a = 16'b1111110111100000;
            14'h6934: o_data_a = 16'b1110110111100000;
            14'h6935: o_data_a = 16'b1111110000010000;
            14'h6936: o_data_a = 16'b0000000000000000;
            14'h6937: o_data_a = 16'b1111110111101000;
            14'h6938: o_data_a = 16'b1110110010100000;
            14'h6939: o_data_a = 16'b1110001100001000;
            14'h693a: o_data_a = 16'b0000000000000000;
            14'h693b: o_data_a = 16'b1111110010101000;
            14'h693c: o_data_a = 16'b1111110000010000;
            14'h693d: o_data_a = 16'b1110110010100000;
            14'h693e: o_data_a = 16'b1111000010001000;
            14'h693f: o_data_a = 16'b0000000000000000;
            14'h6940: o_data_a = 16'b1111110010101000;
            14'h6941: o_data_a = 16'b1111110000010000;
            14'h6942: o_data_a = 16'b0000000000000100;
            14'h6943: o_data_a = 16'b1110001100001000;
            14'h6944: o_data_a = 16'b0000000000000100;
            14'h6945: o_data_a = 16'b1111110000100000;
            14'h6946: o_data_a = 16'b1111110000010000;
            14'h6947: o_data_a = 16'b0000000000000000;
            14'h6948: o_data_a = 16'b1111110111101000;
            14'h6949: o_data_a = 16'b1110110010100000;
            14'h694a: o_data_a = 16'b1110001100001000;
            14'h694b: o_data_a = 16'b0000000000000000;
            14'h694c: o_data_a = 16'b1111110010101000;
            14'h694d: o_data_a = 16'b1111110000010000;
            14'h694e: o_data_a = 16'b0000000000000101;
            14'h694f: o_data_a = 16'b1110001100001000;
            14'h6950: o_data_a = 16'b0000000000000000;
            14'h6951: o_data_a = 16'b1111110010101000;
            14'h6952: o_data_a = 16'b1111110000010000;
            14'h6953: o_data_a = 16'b0000000000000100;
            14'h6954: o_data_a = 16'b1110001100001000;
            14'h6955: o_data_a = 16'b0000000000000101;
            14'h6956: o_data_a = 16'b1111110000010000;
            14'h6957: o_data_a = 16'b0000000000000000;
            14'h6958: o_data_a = 16'b1111110111101000;
            14'h6959: o_data_a = 16'b1110110010100000;
            14'h695a: o_data_a = 16'b1110001100001000;
            14'h695b: o_data_a = 16'b0000000000000000;
            14'h695c: o_data_a = 16'b1111110010101000;
            14'h695d: o_data_a = 16'b1111110000010000;
            14'h695e: o_data_a = 16'b0000000000000100;
            14'h695f: o_data_a = 16'b1111110000100000;
            14'h6960: o_data_a = 16'b1110001100001000;
            14'h6961: o_data_a = 16'b0000000000000011;
            14'h6962: o_data_a = 16'b1111110111100000;
            14'h6963: o_data_a = 16'b1110110111100000;
            14'h6964: o_data_a = 16'b1111110000010000;
            14'h6965: o_data_a = 16'b0000000000000000;
            14'h6966: o_data_a = 16'b1111110111101000;
            14'h6967: o_data_a = 16'b1110110010100000;
            14'h6968: o_data_a = 16'b1110001100001000;
            14'h6969: o_data_a = 16'b0000000000000000;
            14'h696a: o_data_a = 16'b1111110111001000;
            14'h696b: o_data_a = 16'b1111110010100000;
            14'h696c: o_data_a = 16'b1110111111001000;
            14'h696d: o_data_a = 16'b0000000000000000;
            14'h696e: o_data_a = 16'b1111110010101000;
            14'h696f: o_data_a = 16'b1111110000010000;
            14'h6970: o_data_a = 16'b1110110010100000;
            14'h6971: o_data_a = 16'b1111000010001000;
            14'h6972: o_data_a = 16'b0000000000000000;
            14'h6973: o_data_a = 16'b1111110010101000;
            14'h6974: o_data_a = 16'b1111110000010000;
            14'h6975: o_data_a = 16'b0000000000000011;
            14'h6976: o_data_a = 16'b1111110111100000;
            14'h6977: o_data_a = 16'b1110110111100000;
            14'h6978: o_data_a = 16'b1110001100001000;
            14'h6979: o_data_a = 16'b0110100011100110;
            14'h697a: o_data_a = 16'b1110101010000111;
            14'h697b: o_data_a = 16'b0000000000000001;
            14'h697c: o_data_a = 16'b1111110111100000;
            14'h697d: o_data_a = 16'b1110110111100000;
            14'h697e: o_data_a = 16'b1111110000010000;
            14'h697f: o_data_a = 16'b0000000000000000;
            14'h6980: o_data_a = 16'b1111110111101000;
            14'h6981: o_data_a = 16'b1110110010100000;
            14'h6982: o_data_a = 16'b1110001100001000;
            14'h6983: o_data_a = 16'b0000000000000001;
            14'h6984: o_data_a = 16'b1110110000010000;
            14'h6985: o_data_a = 16'b0000000000001101;
            14'h6986: o_data_a = 16'b1110001100001000;
            14'h6987: o_data_a = 16'b0001011011110101;
            14'h6988: o_data_a = 16'b1110110000010000;
            14'h6989: o_data_a = 16'b0000000000001110;
            14'h698a: o_data_a = 16'b1110001100001000;
            14'h698b: o_data_a = 16'b0110100110001111;
            14'h698c: o_data_a = 16'b1110110000010000;
            14'h698d: o_data_a = 16'b0000000001011111;
            14'h698e: o_data_a = 16'b1110101010000111;
            14'h698f: o_data_a = 16'b0000000000000000;
            14'h6990: o_data_a = 16'b1111110010101000;
            14'h6991: o_data_a = 16'b1111110000010000;
            14'h6992: o_data_a = 16'b0000000000000101;
            14'h6993: o_data_a = 16'b1110001100001000;
            14'h6994: o_data_a = 16'b0000000000000000;
            14'h6995: o_data_a = 16'b1111110111001000;
            14'h6996: o_data_a = 16'b1111110010100000;
            14'h6997: o_data_a = 16'b1110101010001000;
            14'h6998: o_data_a = 16'b0000000000110110;
            14'h6999: o_data_a = 16'b1110101010000111;
            14'h699a: o_data_a = 16'b0000000010000000;
            14'h699b: o_data_a = 16'b1110110000010000;
            14'h699c: o_data_a = 16'b0000000000000000;
            14'h699d: o_data_a = 16'b1111110111101000;
            14'h699e: o_data_a = 16'b1110110010100000;
            14'h699f: o_data_a = 16'b1110001100001000;
            14'h69a0: o_data_a = 16'b0000000000110110;
            14'h69a1: o_data_a = 16'b1110101010000111;
            14'h69a2: o_data_a = 16'b0000000010000001;
            14'h69a3: o_data_a = 16'b1110110000010000;
            14'h69a4: o_data_a = 16'b0000000000000000;
            14'h69a5: o_data_a = 16'b1111110111101000;
            14'h69a6: o_data_a = 16'b1110110010100000;
            14'h69a7: o_data_a = 16'b1110001100001000;
            14'h69a8: o_data_a = 16'b0000000000110110;
            14'h69a9: o_data_a = 16'b1110101010000111;
            14'h69aa: o_data_a = 16'b0000000000100010;
            14'h69ab: o_data_a = 16'b1110110000010000;
            14'h69ac: o_data_a = 16'b0000000000000000;
            14'h69ad: o_data_a = 16'b1111110111101000;
            14'h69ae: o_data_a = 16'b1110110010100000;
            14'h69af: o_data_a = 16'b1110001100001000;
            14'h69b0: o_data_a = 16'b0000000000110110;
            14'h69b1: o_data_a = 16'b1110101010000111;
            14'h69b2: o_data_a = 16'b0000000000000000;
            14'h69b3: o_data_a = 16'b1110110000010000;
            14'h69b4: o_data_a = 16'b0000000000001101;
            14'h69b5: o_data_a = 16'b1110001100001000;
            14'h69b6: o_data_a = 16'b0010000100000101;
            14'h69b7: o_data_a = 16'b1110110000010000;
            14'h69b8: o_data_a = 16'b0000000000001110;
            14'h69b9: o_data_a = 16'b1110001100001000;
            14'h69ba: o_data_a = 16'b0110100110111110;
            14'h69bb: o_data_a = 16'b1110110000010000;
            14'h69bc: o_data_a = 16'b0000000001011111;
            14'h69bd: o_data_a = 16'b1110101010000111;
            14'h69be: o_data_a = 16'b0000000000000000;
            14'h69bf: o_data_a = 16'b1111110010101000;
            14'h69c0: o_data_a = 16'b1111110000010000;
            14'h69c1: o_data_a = 16'b0000000000000101;
            14'h69c2: o_data_a = 16'b1110001100001000;
            14'h69c3: o_data_a = 16'b0000000000000000;
            14'h69c4: o_data_a = 16'b1110110000010000;
            14'h69c5: o_data_a = 16'b0000000000001101;
            14'h69c6: o_data_a = 16'b1110001100001000;
            14'h69c7: o_data_a = 16'b0001100101101001;
            14'h69c8: o_data_a = 16'b1110110000010000;
            14'h69c9: o_data_a = 16'b0000000000001110;
            14'h69ca: o_data_a = 16'b1110001100001000;
            14'h69cb: o_data_a = 16'b0110100111001111;
            14'h69cc: o_data_a = 16'b1110110000010000;
            14'h69cd: o_data_a = 16'b0000000001011111;
            14'h69ce: o_data_a = 16'b1110101010000111;
            14'h69cf: o_data_a = 16'b0000000000000000;
            14'h69d0: o_data_a = 16'b1111110010101000;
            14'h69d1: o_data_a = 16'b1111110000010000;
            14'h69d2: o_data_a = 16'b0000000000000101;
            14'h69d3: o_data_a = 16'b1110001100001000;
            14'h69d4: o_data_a = 16'b0000000000000000;
            14'h69d5: o_data_a = 16'b1110110000010000;
            14'h69d6: o_data_a = 16'b0000000000001101;
            14'h69d7: o_data_a = 16'b1110001100001000;
            14'h69d8: o_data_a = 16'b0100111101101001;
            14'h69d9: o_data_a = 16'b1110110000010000;
            14'h69da: o_data_a = 16'b0000000000001110;
            14'h69db: o_data_a = 16'b1110001100001000;
            14'h69dc: o_data_a = 16'b0110100111100000;
            14'h69dd: o_data_a = 16'b1110110000010000;
            14'h69de: o_data_a = 16'b0000000001011111;
            14'h69df: o_data_a = 16'b1110101010000111;
            14'h69e0: o_data_a = 16'b0000000000000000;
            14'h69e1: o_data_a = 16'b1111110010101000;
            14'h69e2: o_data_a = 16'b1111110000010000;
            14'h69e3: o_data_a = 16'b0000000000000101;
            14'h69e4: o_data_a = 16'b1110001100001000;
            14'h69e5: o_data_a = 16'b0000000000000000;
            14'h69e6: o_data_a = 16'b1110110000010000;
            14'h69e7: o_data_a = 16'b0000000000001101;
            14'h69e8: o_data_a = 16'b1110001100001000;
            14'h69e9: o_data_a = 16'b0010011001111110;
            14'h69ea: o_data_a = 16'b1110110000010000;
            14'h69eb: o_data_a = 16'b0000000000001110;
            14'h69ec: o_data_a = 16'b1110001100001000;
            14'h69ed: o_data_a = 16'b0110100111110001;
            14'h69ee: o_data_a = 16'b1110110000010000;
            14'h69ef: o_data_a = 16'b0000000001011111;
            14'h69f0: o_data_a = 16'b1110101010000111;
            14'h69f1: o_data_a = 16'b0000000000000000;
            14'h69f2: o_data_a = 16'b1111110010101000;
            14'h69f3: o_data_a = 16'b1111110000010000;
            14'h69f4: o_data_a = 16'b0000000000000101;
            14'h69f5: o_data_a = 16'b1110001100001000;
            14'h69f6: o_data_a = 16'b0000000000000000;
            14'h69f7: o_data_a = 16'b1110110000010000;
            14'h69f8: o_data_a = 16'b0000000000001101;
            14'h69f9: o_data_a = 16'b1110001100001000;
            14'h69fa: o_data_a = 16'b0001011100011110;
            14'h69fb: o_data_a = 16'b1110110000010000;
            14'h69fc: o_data_a = 16'b0000000000001110;
            14'h69fd: o_data_a = 16'b1110001100001000;
            14'h69fe: o_data_a = 16'b0110101000000010;
            14'h69ff: o_data_a = 16'b1110110000010000;
            14'h6a00: o_data_a = 16'b0000000001011111;
            14'h6a01: o_data_a = 16'b1110101010000111;
            14'h6a02: o_data_a = 16'b0000000000000000;
            14'h6a03: o_data_a = 16'b1111110010101000;
            14'h6a04: o_data_a = 16'b1111110000010000;
            14'h6a05: o_data_a = 16'b0000000000000101;
            14'h6a06: o_data_a = 16'b1110001100001000;
            14'h6a07: o_data_a = 16'b0000000000000000;
            14'h6a08: o_data_a = 16'b1110110000010000;
            14'h6a09: o_data_a = 16'b0000000000001101;
            14'h6a0a: o_data_a = 16'b1110001100001000;
            14'h6a0b: o_data_a = 16'b0000111011111101;
            14'h6a0c: o_data_a = 16'b1110110000010000;
            14'h6a0d: o_data_a = 16'b0000000000001110;
            14'h6a0e: o_data_a = 16'b1110001100001000;
            14'h6a0f: o_data_a = 16'b0110101000010011;
            14'h6a10: o_data_a = 16'b1110110000010000;
            14'h6a11: o_data_a = 16'b0000000001011111;
            14'h6a12: o_data_a = 16'b1110101010000111;
            14'h6a13: o_data_a = 16'b0000000000000000;
            14'h6a14: o_data_a = 16'b1111110010101000;
            14'h6a15: o_data_a = 16'b1111110000010000;
            14'h6a16: o_data_a = 16'b0000000000000101;
            14'h6a17: o_data_a = 16'b1110001100001000;
            14'h6a18: o_data_a = 16'b0000000000000000;
            14'h6a19: o_data_a = 16'b1110110000010000;
            14'h6a1a: o_data_a = 16'b0000000000001101;
            14'h6a1b: o_data_a = 16'b1110001100001000;
            14'h6a1c: o_data_a = 16'b0110101000101001;
            14'h6a1d: o_data_a = 16'b1110110000010000;
            14'h6a1e: o_data_a = 16'b0000000000001110;
            14'h6a1f: o_data_a = 16'b1110001100001000;
            14'h6a20: o_data_a = 16'b0110101000100100;
            14'h6a21: o_data_a = 16'b1110110000010000;
            14'h6a22: o_data_a = 16'b0000000001011111;
            14'h6a23: o_data_a = 16'b1110101010000111;
            14'h6a24: o_data_a = 16'b0000000000000000;
            14'h6a25: o_data_a = 16'b1111110010101000;
            14'h6a26: o_data_a = 16'b1111110000010000;
            14'h6a27: o_data_a = 16'b0000000000000101;
            14'h6a28: o_data_a = 16'b1110001100001000;
            14'h6a29: o_data_a = 16'b0000000000000000;
            14'h6a2a: o_data_a = 16'b1111110111001000;
            14'h6a2b: o_data_a = 16'b1111110010100000;
            14'h6a2c: o_data_a = 16'b1110101010001000;
            14'h6a2d: o_data_a = 16'b0000000000000000;
            14'h6a2e: o_data_a = 16'b1111110010100000;
            14'h6a2f: o_data_a = 16'b1111110001001000;
            14'h6a30: o_data_a = 16'b0000000000000000;
            14'h6a31: o_data_a = 16'b1111110010100000;
            14'h6a32: o_data_a = 16'b1111110001001000;
            14'h6a33: o_data_a = 16'b0000000000000000;
            14'h6a34: o_data_a = 16'b1111110010101000;
            14'h6a35: o_data_a = 16'b1111110000010000;
            14'h6a36: o_data_a = 16'b0110101000111010;
            14'h6a37: o_data_a = 16'b1110001100000101;
            14'h6a38: o_data_a = 16'b0110101000101001;
            14'h6a39: o_data_a = 16'b1110101010000111;
            14'h6a3a: o_data_a = 16'b0000000000000000;
            14'h6a3b: o_data_a = 16'b1111110111101000;
            14'h6a3c: o_data_a = 16'b1110110010100000;
            14'h6a3d: o_data_a = 16'b1110101010001000;
            14'h6a3e: o_data_a = 16'b0000000000000010;
            14'h6a3f: o_data_a = 16'b1111110000100000;
            14'h6a40: o_data_a = 16'b1111110000010000;
            14'h6a41: o_data_a = 16'b0000000000000000;
            14'h6a42: o_data_a = 16'b1111110111101000;
            14'h6a43: o_data_a = 16'b1110110010100000;
            14'h6a44: o_data_a = 16'b1110001100001000;
            14'h6a45: o_data_a = 16'b0000000000000000;
            14'h6a46: o_data_a = 16'b1111110111001000;
            14'h6a47: o_data_a = 16'b1111110010100000;
            14'h6a48: o_data_a = 16'b1110101010001000;
            14'h6a49: o_data_a = 16'b0110101001001101;
            14'h6a4a: o_data_a = 16'b1110110000010000;
            14'h6a4b: o_data_a = 16'b0000000000100110;
            14'h6a4c: o_data_a = 16'b1110101010000111;
            14'h6a4d: o_data_a = 16'b0000000000000000;
            14'h6a4e: o_data_a = 16'b1111110010101000;
            14'h6a4f: o_data_a = 16'b1111110000010000;
            14'h6a50: o_data_a = 16'b0110101001010100;
            14'h6a51: o_data_a = 16'b1110001100000101;
            14'h6a52: o_data_a = 16'b0110101001101001;
            14'h6a53: o_data_a = 16'b1110101010000111;
            14'h6a54: o_data_a = 16'b0000000000000000;
            14'h6a55: o_data_a = 16'b1111110111001000;
            14'h6a56: o_data_a = 16'b1111110010100000;
            14'h6a57: o_data_a = 16'b1110111111001000;
            14'h6a58: o_data_a = 16'b0000000000000001;
            14'h6a59: o_data_a = 16'b1110110000010000;
            14'h6a5a: o_data_a = 16'b0000000000001101;
            14'h6a5b: o_data_a = 16'b1110001100001000;
            14'h6a5c: o_data_a = 16'b0110101011011001;
            14'h6a5d: o_data_a = 16'b1110110000010000;
            14'h6a5e: o_data_a = 16'b0000000000001110;
            14'h6a5f: o_data_a = 16'b1110001100001000;
            14'h6a60: o_data_a = 16'b0110101001100100;
            14'h6a61: o_data_a = 16'b1110110000010000;
            14'h6a62: o_data_a = 16'b0000000001011111;
            14'h6a63: o_data_a = 16'b1110101010000111;
            14'h6a64: o_data_a = 16'b0000000000000000;
            14'h6a65: o_data_a = 16'b1111110010101000;
            14'h6a66: o_data_a = 16'b1111110000010000;
            14'h6a67: o_data_a = 16'b0000000000000101;
            14'h6a68: o_data_a = 16'b1110001100001000;
            14'h6a69: o_data_a = 16'b0000000000000010;
            14'h6a6a: o_data_a = 16'b1111110000100000;
            14'h6a6b: o_data_a = 16'b1111110000010000;
            14'h6a6c: o_data_a = 16'b0000000000000000;
            14'h6a6d: o_data_a = 16'b1111110111101000;
            14'h6a6e: o_data_a = 16'b1110110010100000;
            14'h6a6f: o_data_a = 16'b1110001100001000;
            14'h6a70: o_data_a = 16'b0000000000000000;
            14'h6a71: o_data_a = 16'b1111110111001000;
            14'h6a72: o_data_a = 16'b1111110010100000;
            14'h6a73: o_data_a = 16'b1110101010001000;
            14'h6a74: o_data_a = 16'b0110101001111000;
            14'h6a75: o_data_a = 16'b1110110000010000;
            14'h6a76: o_data_a = 16'b0000000000010110;
            14'h6a77: o_data_a = 16'b1110101010000111;
            14'h6a78: o_data_a = 16'b0000000000000000;
            14'h6a79: o_data_a = 16'b1111110010100000;
            14'h6a7a: o_data_a = 16'b1111110001001000;
            14'h6a7b: o_data_a = 16'b0000000000000000;
            14'h6a7c: o_data_a = 16'b1111110010101000;
            14'h6a7d: o_data_a = 16'b1111110000010000;
            14'h6a7e: o_data_a = 16'b0110101011010011;
            14'h6a7f: o_data_a = 16'b1110001100000101;
            14'h6a80: o_data_a = 16'b0000000000110010;
            14'h6a81: o_data_a = 16'b1110110000010000;
            14'h6a82: o_data_a = 16'b0000000000000000;
            14'h6a83: o_data_a = 16'b1111110111101000;
            14'h6a84: o_data_a = 16'b1110110010100000;
            14'h6a85: o_data_a = 16'b1110001100001000;
            14'h6a86: o_data_a = 16'b0000000000000000;
            14'h6a87: o_data_a = 16'b1111110010101000;
            14'h6a88: o_data_a = 16'b1111110000010000;
            14'h6a89: o_data_a = 16'b0000000000000001;
            14'h6a8a: o_data_a = 16'b1111110000100000;
            14'h6a8b: o_data_a = 16'b1110001100001000;
            14'h6a8c: o_data_a = 16'b0000000000000001;
            14'h6a8d: o_data_a = 16'b1111110000100000;
            14'h6a8e: o_data_a = 16'b1111110000010000;
            14'h6a8f: o_data_a = 16'b0000000000000000;
            14'h6a90: o_data_a = 16'b1111110111101000;
            14'h6a91: o_data_a = 16'b1110110010100000;
            14'h6a92: o_data_a = 16'b1110001100001000;
            14'h6a93: o_data_a = 16'b0000000000000000;
            14'h6a94: o_data_a = 16'b1111110111001000;
            14'h6a95: o_data_a = 16'b1111110010100000;
            14'h6a96: o_data_a = 16'b1110101010001000;
            14'h6a97: o_data_a = 16'b0110101010011011;
            14'h6a98: o_data_a = 16'b1110110000010000;
            14'h6a99: o_data_a = 16'b0000000000010110;
            14'h6a9a: o_data_a = 16'b1110101010000111;
            14'h6a9b: o_data_a = 16'b0000000000000000;
            14'h6a9c: o_data_a = 16'b1111110010100000;
            14'h6a9d: o_data_a = 16'b1111110001001000;
            14'h6a9e: o_data_a = 16'b0000000000000000;
            14'h6a9f: o_data_a = 16'b1111110010101000;
            14'h6aa0: o_data_a = 16'b1111110000010000;
            14'h6aa1: o_data_a = 16'b0110101010111011;
            14'h6aa2: o_data_a = 16'b1110001100000101;
            14'h6aa3: o_data_a = 16'b0000000000000001;
            14'h6aa4: o_data_a = 16'b1111110000100000;
            14'h6aa5: o_data_a = 16'b1111110000010000;
            14'h6aa6: o_data_a = 16'b0000000000000000;
            14'h6aa7: o_data_a = 16'b1111110111101000;
            14'h6aa8: o_data_a = 16'b1110110010100000;
            14'h6aa9: o_data_a = 16'b1110001100001000;
            14'h6aaa: o_data_a = 16'b0000000000000000;
            14'h6aab: o_data_a = 16'b1111110111001000;
            14'h6aac: o_data_a = 16'b1111110010100000;
            14'h6aad: o_data_a = 16'b1110111111001000;
            14'h6aae: o_data_a = 16'b0000000000000000;
            14'h6aaf: o_data_a = 16'b1111110010101000;
            14'h6ab0: o_data_a = 16'b1111110000010000;
            14'h6ab1: o_data_a = 16'b1110110010100000;
            14'h6ab2: o_data_a = 16'b1111000111001000;
            14'h6ab3: o_data_a = 16'b0000000000000000;
            14'h6ab4: o_data_a = 16'b1111110010101000;
            14'h6ab5: o_data_a = 16'b1111110000010000;
            14'h6ab6: o_data_a = 16'b0000000000000001;
            14'h6ab7: o_data_a = 16'b1111110000100000;
            14'h6ab8: o_data_a = 16'b1110001100001000;
            14'h6ab9: o_data_a = 16'b0110101010001100;
            14'h6aba: o_data_a = 16'b1110101010000111;
            14'h6abb: o_data_a = 16'b0000000000000010;
            14'h6abc: o_data_a = 16'b1111110000100000;
            14'h6abd: o_data_a = 16'b1111110000010000;
            14'h6abe: o_data_a = 16'b0000000000000000;
            14'h6abf: o_data_a = 16'b1111110111101000;
            14'h6ac0: o_data_a = 16'b1110110010100000;
            14'h6ac1: o_data_a = 16'b1110001100001000;
            14'h6ac2: o_data_a = 16'b0000000000000000;
            14'h6ac3: o_data_a = 16'b1111110111001000;
            14'h6ac4: o_data_a = 16'b1111110010100000;
            14'h6ac5: o_data_a = 16'b1110111111001000;
            14'h6ac6: o_data_a = 16'b0000000000000000;
            14'h6ac7: o_data_a = 16'b1111110010101000;
            14'h6ac8: o_data_a = 16'b1111110000010000;
            14'h6ac9: o_data_a = 16'b1110110010100000;
            14'h6aca: o_data_a = 16'b1111000111001000;
            14'h6acb: o_data_a = 16'b0000000000000000;
            14'h6acc: o_data_a = 16'b1111110010101000;
            14'h6acd: o_data_a = 16'b1111110000010000;
            14'h6ace: o_data_a = 16'b0000000000000010;
            14'h6acf: o_data_a = 16'b1111110000100000;
            14'h6ad0: o_data_a = 16'b1110001100001000;
            14'h6ad1: o_data_a = 16'b0110101001101001;
            14'h6ad2: o_data_a = 16'b1110101010000111;
            14'h6ad3: o_data_a = 16'b0000000000000000;
            14'h6ad4: o_data_a = 16'b1111110111001000;
            14'h6ad5: o_data_a = 16'b1111110010100000;
            14'h6ad6: o_data_a = 16'b1110101010001000;
            14'h6ad7: o_data_a = 16'b0000000000110110;
            14'h6ad8: o_data_a = 16'b1110101010000111;
            14'h6ad9: o_data_a = 16'b0000000000000011;
            14'h6ada: o_data_a = 16'b1110110000010000;
            14'h6adb: o_data_a = 16'b0000000000000000;
            14'h6adc: o_data_a = 16'b1111110111101000;
            14'h6add: o_data_a = 16'b1110110010100000;
            14'h6ade: o_data_a = 16'b1110001100001000;
            14'h6adf: o_data_a = 16'b0000000000000001;
            14'h6ae0: o_data_a = 16'b1110110000010000;
            14'h6ae1: o_data_a = 16'b0000000000001101;
            14'h6ae2: o_data_a = 16'b1110001100001000;
            14'h6ae3: o_data_a = 16'b0110001000010001;
            14'h6ae4: o_data_a = 16'b1110110000010000;
            14'h6ae5: o_data_a = 16'b0000000000001110;
            14'h6ae6: o_data_a = 16'b1110001100001000;
            14'h6ae7: o_data_a = 16'b0110101011101011;
            14'h6ae8: o_data_a = 16'b1110110000010000;
            14'h6ae9: o_data_a = 16'b0000000001011111;
            14'h6aea: o_data_a = 16'b1110101010000111;
            14'h6aeb: o_data_a = 16'b0000000001000101;
            14'h6aec: o_data_a = 16'b1110110000010000;
            14'h6aed: o_data_a = 16'b0000000000000000;
            14'h6aee: o_data_a = 16'b1111110111101000;
            14'h6aef: o_data_a = 16'b1110110010100000;
            14'h6af0: o_data_a = 16'b1110001100001000;
            14'h6af1: o_data_a = 16'b0000000000000010;
            14'h6af2: o_data_a = 16'b1110110000010000;
            14'h6af3: o_data_a = 16'b0000000000001101;
            14'h6af4: o_data_a = 16'b1110001100001000;
            14'h6af5: o_data_a = 16'b0110010000111011;
            14'h6af6: o_data_a = 16'b1110110000010000;
            14'h6af7: o_data_a = 16'b0000000000001110;
            14'h6af8: o_data_a = 16'b1110001100001000;
            14'h6af9: o_data_a = 16'b0110101011111101;
            14'h6afa: o_data_a = 16'b1110110000010000;
            14'h6afb: o_data_a = 16'b0000000001011111;
            14'h6afc: o_data_a = 16'b1110101010000111;
            14'h6afd: o_data_a = 16'b0000000001010010;
            14'h6afe: o_data_a = 16'b1110110000010000;
            14'h6aff: o_data_a = 16'b0000000000000000;
            14'h6b00: o_data_a = 16'b1111110111101000;
            14'h6b01: o_data_a = 16'b1110110010100000;
            14'h6b02: o_data_a = 16'b1110001100001000;
            14'h6b03: o_data_a = 16'b0000000000000010;
            14'h6b04: o_data_a = 16'b1110110000010000;
            14'h6b05: o_data_a = 16'b0000000000001101;
            14'h6b06: o_data_a = 16'b1110001100001000;
            14'h6b07: o_data_a = 16'b0110010000111011;
            14'h6b08: o_data_a = 16'b1110110000010000;
            14'h6b09: o_data_a = 16'b0000000000001110;
            14'h6b0a: o_data_a = 16'b1110001100001000;
            14'h6b0b: o_data_a = 16'b0110101100001111;
            14'h6b0c: o_data_a = 16'b1110110000010000;
            14'h6b0d: o_data_a = 16'b0000000001011111;
            14'h6b0e: o_data_a = 16'b1110101010000111;
            14'h6b0f: o_data_a = 16'b0000000001010010;
            14'h6b10: o_data_a = 16'b1110110000010000;
            14'h6b11: o_data_a = 16'b0000000000000000;
            14'h6b12: o_data_a = 16'b1111110111101000;
            14'h6b13: o_data_a = 16'b1110110010100000;
            14'h6b14: o_data_a = 16'b1110001100001000;
            14'h6b15: o_data_a = 16'b0000000000000010;
            14'h6b16: o_data_a = 16'b1110110000010000;
            14'h6b17: o_data_a = 16'b0000000000001101;
            14'h6b18: o_data_a = 16'b1110001100001000;
            14'h6b19: o_data_a = 16'b0110010000111011;
            14'h6b1a: o_data_a = 16'b1110110000010000;
            14'h6b1b: o_data_a = 16'b0000000000001110;
            14'h6b1c: o_data_a = 16'b1110001100001000;
            14'h6b1d: o_data_a = 16'b0110101100100001;
            14'h6b1e: o_data_a = 16'b1110110000010000;
            14'h6b1f: o_data_a = 16'b0000000001011111;
            14'h6b20: o_data_a = 16'b1110101010000111;
            14'h6b21: o_data_a = 16'b0000000000000001;
            14'h6b22: o_data_a = 16'b1110110000010000;
            14'h6b23: o_data_a = 16'b0000000000001101;
            14'h6b24: o_data_a = 16'b1110001100001000;
            14'h6b25: o_data_a = 16'b0100110110001010;
            14'h6b26: o_data_a = 16'b1110110000010000;
            14'h6b27: o_data_a = 16'b0000000000001110;
            14'h6b28: o_data_a = 16'b1110001100001000;
            14'h6b29: o_data_a = 16'b0110101100101101;
            14'h6b2a: o_data_a = 16'b1110110000010000;
            14'h6b2b: o_data_a = 16'b0000000001011111;
            14'h6b2c: o_data_a = 16'b1110101010000111;
            14'h6b2d: o_data_a = 16'b0000000000000000;
            14'h6b2e: o_data_a = 16'b1111110010101000;
            14'h6b2f: o_data_a = 16'b1111110000010000;
            14'h6b30: o_data_a = 16'b0000000000000101;
            14'h6b31: o_data_a = 16'b1110001100001000;
            14'h6b32: o_data_a = 16'b0000000000000010;
            14'h6b33: o_data_a = 16'b1111110000100000;
            14'h6b34: o_data_a = 16'b1111110000010000;
            14'h6b35: o_data_a = 16'b0000000000000000;
            14'h6b36: o_data_a = 16'b1111110111101000;
            14'h6b37: o_data_a = 16'b1110110010100000;
            14'h6b38: o_data_a = 16'b1110001100001000;
            14'h6b39: o_data_a = 16'b0000000000000001;
            14'h6b3a: o_data_a = 16'b1110110000010000;
            14'h6b3b: o_data_a = 16'b0000000000001101;
            14'h6b3c: o_data_a = 16'b1110001100001000;
            14'h6b3d: o_data_a = 16'b0100111000001101;
            14'h6b3e: o_data_a = 16'b1110110000010000;
            14'h6b3f: o_data_a = 16'b0000000000001110;
            14'h6b40: o_data_a = 16'b1110001100001000;
            14'h6b41: o_data_a = 16'b0110101101000101;
            14'h6b42: o_data_a = 16'b1110110000010000;
            14'h6b43: o_data_a = 16'b0000000001011111;
            14'h6b44: o_data_a = 16'b1110101010000111;
            14'h6b45: o_data_a = 16'b0000000000000000;
            14'h6b46: o_data_a = 16'b1111110010101000;
            14'h6b47: o_data_a = 16'b1111110000010000;
            14'h6b48: o_data_a = 16'b0000000000000101;
            14'h6b49: o_data_a = 16'b1110001100001000;
            14'h6b4a: o_data_a = 16'b0000000000000000;
            14'h6b4b: o_data_a = 16'b1110110000010000;
            14'h6b4c: o_data_a = 16'b0000000000001101;
            14'h6b4d: o_data_a = 16'b1110001100001000;
            14'h6b4e: o_data_a = 16'b0110101000101001;
            14'h6b4f: o_data_a = 16'b1110110000010000;
            14'h6b50: o_data_a = 16'b0000000000001110;
            14'h6b51: o_data_a = 16'b1110001100001000;
            14'h6b52: o_data_a = 16'b0110101101010110;
            14'h6b53: o_data_a = 16'b1110110000010000;
            14'h6b54: o_data_a = 16'b0000000001011111;
            14'h6b55: o_data_a = 16'b1110101010000111;
            14'h6b56: o_data_a = 16'b0000000000000000;
            14'h6b57: o_data_a = 16'b1111110010101000;
            14'h6b58: o_data_a = 16'b1111110000010000;
            14'h6b59: o_data_a = 16'b0000000000000101;
            14'h6b5a: o_data_a = 16'b1110001100001000;
            default: o_data_a = 16'b0000000000000000;
       endcase
   end 

endmodule
